

module i1s11
(
  input DIN,
  input DIN_t,
  output Q,
  output Q_t
);

  assign Q = ~DIN;
  assign Q_t = DIN_t;

endmodule



module and2s1
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  output Q,
  output Q_t
);

  assign Q = DIN1 & DIN2;
  assign Q_t = DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1);

endmodule



module or4s1
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  input DIN3,
  input DIN3_t,
  input DIN4,
  input DIN4_t,
  output Q,
  output Q_t
);

  assign Q = DIN1 | DIN2 | DIN3 | DIN4;
  assign Q_t = ((DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1)) & DIN3_t | ((DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1)) & ~DIN3 | DIN3_t & ~(DIN1 | DIN2))) & DIN4_t | (((DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1)) & DIN3_t | ((DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1)) & ~DIN3 | DIN3_t & ~(DIN1 | DIN2))) & ~DIN4 | DIN4_t & ~(DIN1 | DIN2 | DIN3));

endmodule



module i1s3
(
  input DIN,
  input DIN_t,
  output Q,
  output Q_t
);

  assign Q = ~DIN;
  assign Q_t = DIN_t;

endmodule



module or3s1
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  input DIN3,
  input DIN3_t,
  output Q,
  output Q_t
);

  assign Q = DIN1 | DIN2 | DIN3;
  assign Q_t = (DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1)) & DIN3_t | ((DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1)) & ~DIN3 | DIN3_t & ~(DIN1 | DIN2));

endmodule



module i1s1
(
  input DIN,
  input DIN_t,
  output Q,
  output Q_t
);

  assign Q = ~DIN;
  assign Q_t = DIN_t;

endmodule



module i1s12
(
  input DIN,
  input DIN_t,
  output Q,
  output Q_t
);

  assign Q = ~DIN;
  assign Q_t = DIN_t;

endmodule



module nnd4s1
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  input DIN3,
  input DIN3_t,
  input DIN4,
  input DIN4_t,
  output Q,
  output Q_t
);

  assign Q = ~(DIN1 & DIN2 & DIN3 & DIN4);
  assign Q_t = ((DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1)) & DIN3_t | ((DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1)) & DIN3 | DIN3_t & (DIN1 & DIN2))) & DIN4_t | (((DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1)) & DIN3_t | ((DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1)) & DIN3 | DIN3_t & (DIN1 & DIN2))) & DIN4 | DIN4_t & (DIN1 & DIN2 & DIN3));

endmodule



module and2s3
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  output Q,
  output Q_t
);

  assign Q = DIN1 & DIN2;
  assign Q_t = DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1);

endmodule



module nnd2s3
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  output Q,
  output Q_t
);

  assign Q = ~(DIN1 & DIN2);
  assign Q_t = DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1);

endmodule



module ib1s9
(
  input DIN,
  input DIN_t,
  output Q,
  output Q_t
);

  assign Q = DIN;
  assign Q_t = DIN_t;

endmodule



module xor2s1
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  output Q,
  output Q_t
);

  assign Q = DIN1 ^ DIN2;
  assign Q_t = DIN1_t | DIN2_t;

endmodule



module xnr2s3
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  output Q,
  output Q_t
);

  assign Q = ~(DIN1 ^ DIN2);
  assign Q_t = DIN1_t | DIN2_t;

endmodule



module xor2s3
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  output Q,
  output Q_t
);

  assign Q = DIN1 ^ DIN2;
  assign Q_t = DIN1_t | DIN2_t;

endmodule



module sdffs1
(
  input DIN,
  input DIN_t,
  input SDIN,
  input SDIN_t,
  input SSEL,
  input SSEL_t,
  input CLK,
  input CLK_t,
  output reg Q,
  output reg Q_t,
  output QN,
  output QN_t
);


  always @(posedge CLK) begin
    if(SSEL) Q <= SDIN; 
    else Q <= DIN;
  end

  assign QN = ~Q;
  assign QN_t = Q_t;

endmodule



module nor2s3
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  output Q,
  output Q_t
);

  assign Q = ~(DIN1 | DIN2);
  assign Q_t = DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1);

endmodule



module nor4s1
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  input DIN3,
  input DIN3_t,
  input DIN4,
  input DIN4_t,
  output Q,
  output Q_t
);

  assign Q = ~(DIN1 | DIN2 | DIN3 | DIN4);
  assign Q_t = ((DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1)) & DIN3_t | ((DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1)) & ~DIN3 | DIN3_t & ~(DIN1 | DIN2))) & DIN4_t | (((DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1)) & DIN3_t | ((DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1)) & ~DIN3 | DIN3_t & ~(DIN1 | DIN2))) & ~DIN4 | DIN4_t & ~(DIN1 | DIN2 | DIN3));

endmodule



module and3s3
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  input DIN3,
  input DIN3_t,
  output Q,
  output Q_t
);

  assign Q = DIN1 & DIN2 & DIN3;
  assign Q_t = (DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1)) & DIN3_t | ((DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1)) & DIN3 | DIN3_t & (DIN1 & DIN2));

endmodule



module nnd4s2
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  input DIN3,
  input DIN3_t,
  input DIN4,
  input DIN4_t,
  output Q,
  output Q_t
);

  assign Q = ~(DIN1 & DIN2 & DIN3 & DIN4);
  assign Q_t = ((DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1)) & DIN3_t | ((DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1)) & DIN3 | DIN3_t & (DIN1 & DIN2))) & DIN4_t | (((DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1)) & DIN3_t | ((DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1)) & DIN3 | DIN3_t & (DIN1 & DIN2))) & DIN4 | DIN4_t & (DIN1 & DIN2 & DIN3));

endmodule



module nnd2s1
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  output Q,
  output Q_t
);

  assign Q = ~(DIN1 & DIN2);
  assign Q_t = DIN1_t & DIN2_t | (DIN1_t & DIN2 | DIN2_t & DIN1);

endmodule



module nor2s1
(
  input DIN1,
  input DIN1_t,
  input DIN2,
  input DIN2_t,
  output Q,
  output Q_t
);

  assign Q = ~(DIN1 | DIN2);
  assign Q_t = DIN1_t & DIN2_t | (DIN1_t & ~DIN2 | DIN2_t & ~DIN1);

endmodule



module s35932
(
  CK,
  CRC_OUT_1_0,
  CRC_OUT_1_1,
  CRC_OUT_1_10,
  CRC_OUT_1_11,
  CRC_OUT_1_12,
  CRC_OUT_1_13,
  CRC_OUT_1_14,
  CRC_OUT_1_15,
  CRC_OUT_1_16,
  CRC_OUT_1_17,
  CRC_OUT_1_18,
  CRC_OUT_1_19,
  CRC_OUT_1_2,
  CRC_OUT_1_20,
  CRC_OUT_1_21,
  CRC_OUT_1_22,
  CRC_OUT_1_23,
  CRC_OUT_1_24,
  CRC_OUT_1_25,
  CRC_OUT_1_26,
  CRC_OUT_1_27,
  CRC_OUT_1_28,
  CRC_OUT_1_29,
  CRC_OUT_1_3,
  CRC_OUT_1_30,
  CRC_OUT_1_31,
  CRC_OUT_1_4,
  CRC_OUT_1_5,
  CRC_OUT_1_6,
  CRC_OUT_1_7,
  CRC_OUT_1_8,
  CRC_OUT_1_9,
  CRC_OUT_2_0,
  CRC_OUT_2_1,
  CRC_OUT_2_10,
  CRC_OUT_2_11,
  CRC_OUT_2_12,
  CRC_OUT_2_13,
  CRC_OUT_2_14,
  CRC_OUT_2_15,
  CRC_OUT_2_16,
  CRC_OUT_2_17,
  CRC_OUT_2_18,
  CRC_OUT_2_19,
  CRC_OUT_2_2,
  CRC_OUT_2_20,
  CRC_OUT_2_21,
  CRC_OUT_2_22,
  CRC_OUT_2_23,
  CRC_OUT_2_24,
  CRC_OUT_2_25,
  CRC_OUT_2_26,
  CRC_OUT_2_27,
  CRC_OUT_2_28,
  CRC_OUT_2_29,
  CRC_OUT_2_3,
  CRC_OUT_2_30,
  CRC_OUT_2_31,
  CRC_OUT_2_4,
  CRC_OUT_2_5,
  CRC_OUT_2_6,
  CRC_OUT_2_7,
  CRC_OUT_2_8,
  CRC_OUT_2_9,
  CRC_OUT_3_0,
  CRC_OUT_3_1,
  CRC_OUT_3_10,
  CRC_OUT_3_11,
  CRC_OUT_3_12,
  CRC_OUT_3_13,
  CRC_OUT_3_14,
  CRC_OUT_3_15,
  CRC_OUT_3_16,
  CRC_OUT_3_17,
  CRC_OUT_3_18,
  CRC_OUT_3_19,
  CRC_OUT_3_2,
  CRC_OUT_3_20,
  CRC_OUT_3_21,
  CRC_OUT_3_22,
  CRC_OUT_3_23,
  CRC_OUT_3_24,
  CRC_OUT_3_25,
  CRC_OUT_3_26,
  CRC_OUT_3_27,
  CRC_OUT_3_28,
  CRC_OUT_3_29,
  CRC_OUT_3_3,
  CRC_OUT_3_30,
  CRC_OUT_3_31,
  CRC_OUT_3_4,
  CRC_OUT_3_5,
  CRC_OUT_3_6,
  CRC_OUT_3_7,
  CRC_OUT_3_8,
  CRC_OUT_3_9,
  CRC_OUT_4_0,
  CRC_OUT_4_1,
  CRC_OUT_4_10,
  CRC_OUT_4_11,
  CRC_OUT_4_12,
  CRC_OUT_4_13,
  CRC_OUT_4_14,
  CRC_OUT_4_15,
  CRC_OUT_4_16,
  CRC_OUT_4_17,
  CRC_OUT_4_18,
  CRC_OUT_4_19,
  CRC_OUT_4_2,
  CRC_OUT_4_20,
  CRC_OUT_4_21,
  CRC_OUT_4_22,
  CRC_OUT_4_23,
  CRC_OUT_4_24,
  CRC_OUT_4_25,
  CRC_OUT_4_26,
  CRC_OUT_4_27,
  CRC_OUT_4_28,
  CRC_OUT_4_29,
  CRC_OUT_4_3,
  CRC_OUT_4_30,
  CRC_OUT_4_31,
  CRC_OUT_4_4,
  CRC_OUT_4_5,
  CRC_OUT_4_6,
  CRC_OUT_4_7,
  CRC_OUT_4_8,
  CRC_OUT_4_9,
  CRC_OUT_5_0,
  CRC_OUT_5_1,
  CRC_OUT_5_10,
  CRC_OUT_5_11,
  CRC_OUT_5_12,
  CRC_OUT_5_13,
  CRC_OUT_5_14,
  CRC_OUT_5_15,
  CRC_OUT_5_16,
  CRC_OUT_5_17,
  CRC_OUT_5_18,
  CRC_OUT_5_19,
  CRC_OUT_5_2,
  CRC_OUT_5_20,
  CRC_OUT_5_21,
  CRC_OUT_5_22,
  CRC_OUT_5_23,
  CRC_OUT_5_24,
  CRC_OUT_5_25,
  CRC_OUT_5_26,
  CRC_OUT_5_27,
  CRC_OUT_5_28,
  CRC_OUT_5_29,
  CRC_OUT_5_3,
  CRC_OUT_5_30,
  CRC_OUT_5_31,
  CRC_OUT_5_4,
  CRC_OUT_5_5,
  CRC_OUT_5_6,
  CRC_OUT_5_7,
  CRC_OUT_5_8,
  CRC_OUT_5_9,
  CRC_OUT_6_0,
  CRC_OUT_6_1,
  CRC_OUT_6_10,
  CRC_OUT_6_11,
  CRC_OUT_6_12,
  CRC_OUT_6_13,
  CRC_OUT_6_14,
  CRC_OUT_6_15,
  CRC_OUT_6_16,
  CRC_OUT_6_17,
  CRC_OUT_6_18,
  CRC_OUT_6_19,
  CRC_OUT_6_2,
  CRC_OUT_6_20,
  CRC_OUT_6_21,
  CRC_OUT_6_22,
  CRC_OUT_6_23,
  CRC_OUT_6_24,
  CRC_OUT_6_25,
  CRC_OUT_6_26,
  CRC_OUT_6_27,
  CRC_OUT_6_28,
  CRC_OUT_6_29,
  CRC_OUT_6_3,
  CRC_OUT_6_30,
  CRC_OUT_6_31,
  CRC_OUT_6_4,
  CRC_OUT_6_5,
  CRC_OUT_6_6,
  CRC_OUT_6_7,
  CRC_OUT_6_8,
  CRC_OUT_6_9,
  CRC_OUT_7_0,
  CRC_OUT_7_1,
  CRC_OUT_7_10,
  CRC_OUT_7_11,
  CRC_OUT_7_12,
  CRC_OUT_7_13,
  CRC_OUT_7_14,
  CRC_OUT_7_15,
  CRC_OUT_7_16,
  CRC_OUT_7_17,
  CRC_OUT_7_18,
  CRC_OUT_7_19,
  CRC_OUT_7_2,
  CRC_OUT_7_20,
  CRC_OUT_7_21,
  CRC_OUT_7_22,
  CRC_OUT_7_23,
  CRC_OUT_7_24,
  CRC_OUT_7_25,
  CRC_OUT_7_26,
  CRC_OUT_7_27,
  CRC_OUT_7_28,
  CRC_OUT_7_29,
  CRC_OUT_7_3,
  CRC_OUT_7_30,
  CRC_OUT_7_31,
  CRC_OUT_7_4,
  CRC_OUT_7_5,
  CRC_OUT_7_6,
  CRC_OUT_7_7,
  CRC_OUT_7_8,
  CRC_OUT_7_9,
  CRC_OUT_8_0,
  CRC_OUT_8_1,
  CRC_OUT_8_10,
  CRC_OUT_8_11,
  CRC_OUT_8_12,
  CRC_OUT_8_13,
  CRC_OUT_8_14,
  CRC_OUT_8_15,
  CRC_OUT_8_16,
  CRC_OUT_8_17,
  CRC_OUT_8_18,
  CRC_OUT_8_19,
  CRC_OUT_8_2,
  CRC_OUT_8_20,
  CRC_OUT_8_21,
  CRC_OUT_8_22,
  CRC_OUT_8_23,
  CRC_OUT_8_24,
  CRC_OUT_8_25,
  CRC_OUT_8_26,
  CRC_OUT_8_27,
  CRC_OUT_8_28,
  CRC_OUT_8_29,
  CRC_OUT_8_3,
  CRC_OUT_8_30,
  CRC_OUT_8_31,
  CRC_OUT_8_4,
  CRC_OUT_8_5,
  CRC_OUT_8_6,
  CRC_OUT_8_7,
  CRC_OUT_8_8,
  CRC_OUT_8_9,
  CRC_OUT_9_0,
  CRC_OUT_9_1,
  CRC_OUT_9_10,
  CRC_OUT_9_11,
  CRC_OUT_9_12,
  CRC_OUT_9_13,
  CRC_OUT_9_14,
  CRC_OUT_9_15,
  CRC_OUT_9_16,
  CRC_OUT_9_17,
  CRC_OUT_9_18,
  CRC_OUT_9_19,
  CRC_OUT_9_2,
  CRC_OUT_9_20,
  CRC_OUT_9_21,
  CRC_OUT_9_22,
  CRC_OUT_9_23,
  CRC_OUT_9_24,
  CRC_OUT_9_25,
  CRC_OUT_9_26,
  CRC_OUT_9_27,
  CRC_OUT_9_28,
  CRC_OUT_9_29,
  CRC_OUT_9_3,
  CRC_OUT_9_30,
  CRC_OUT_9_31,
  CRC_OUT_9_4,
  CRC_OUT_9_5,
  CRC_OUT_9_6,
  CRC_OUT_9_7,
  CRC_OUT_9_8,
  CRC_OUT_9_9,
  DATA_0_0,
  DATA_0_1,
  DATA_0_10,
  DATA_0_11,
  DATA_0_12,
  DATA_0_13,
  DATA_0_14,
  DATA_0_15,
  DATA_0_16,
  DATA_0_17,
  DATA_0_18,
  DATA_0_19,
  DATA_0_2,
  DATA_0_20,
  DATA_0_21,
  DATA_0_22,
  DATA_0_23,
  DATA_0_24,
  DATA_0_25,
  DATA_0_26,
  DATA_0_27,
  DATA_0_28,
  DATA_0_29,
  DATA_0_3,
  DATA_0_30,
  DATA_0_31,
  DATA_0_4,
  DATA_0_5,
  DATA_0_6,
  DATA_0_7,
  DATA_0_8,
  DATA_0_9,
  DATA_9_0,
  DATA_9_1,
  DATA_9_10,
  DATA_9_11,
  DATA_9_12,
  DATA_9_13,
  DATA_9_14,
  DATA_9_15,
  DATA_9_16,
  DATA_9_17,
  DATA_9_18,
  DATA_9_19,
  DATA_9_2,
  DATA_9_20,
  DATA_9_21,
  DATA_9_22,
  DATA_9_23,
  DATA_9_24,
  DATA_9_25,
  DATA_9_26,
  DATA_9_27,
  DATA_9_28,
  DATA_9_29,
  DATA_9_3,
  DATA_9_30,
  DATA_9_31,
  DATA_9_4,
  DATA_9_5,
  DATA_9_6,
  DATA_9_7,
  DATA_9_8,
  DATA_9_9,
  RESET,
  TM0,
  TM1,
  test_se,
  test_si,
  test_so
);

  input CK;input DATA_0_0;input DATA_0_1;input DATA_0_10;input DATA_0_11;input DATA_0_12;input DATA_0_13;input DATA_0_14;input DATA_0_15;input DATA_0_16;input DATA_0_17;input DATA_0_18;input DATA_0_19;input DATA_0_2;input DATA_0_20;input DATA_0_21;input DATA_0_22;input DATA_0_23;input DATA_0_24;input DATA_0_25;input DATA_0_26;input DATA_0_27;input DATA_0_28;input DATA_0_29;input DATA_0_3;input DATA_0_30;input DATA_0_31;input DATA_0_4;input DATA_0_5;input DATA_0_6;input DATA_0_7;input DATA_0_8;input DATA_0_9;input RESET;input TM0;input TM1;input test_se;input test_si;
  output CRC_OUT_1_0;output CRC_OUT_1_1;output CRC_OUT_1_10;output CRC_OUT_1_11;output CRC_OUT_1_12;output CRC_OUT_1_13;output CRC_OUT_1_14;output CRC_OUT_1_15;output CRC_OUT_1_16;output CRC_OUT_1_17;output CRC_OUT_1_18;output CRC_OUT_1_19;output CRC_OUT_1_2;output CRC_OUT_1_20;output CRC_OUT_1_21;output CRC_OUT_1_22;output CRC_OUT_1_23;output CRC_OUT_1_24;output CRC_OUT_1_25;output CRC_OUT_1_26;output CRC_OUT_1_27;output CRC_OUT_1_28;output CRC_OUT_1_29;output CRC_OUT_1_3;output CRC_OUT_1_30;output CRC_OUT_1_31;output CRC_OUT_1_4;output CRC_OUT_1_5;output CRC_OUT_1_6;output CRC_OUT_1_7;output CRC_OUT_1_8;output CRC_OUT_1_9;output CRC_OUT_2_0;output CRC_OUT_2_1;output CRC_OUT_2_10;output CRC_OUT_2_11;output CRC_OUT_2_12;output CRC_OUT_2_13;output CRC_OUT_2_14;output CRC_OUT_2_15;output CRC_OUT_2_16;output CRC_OUT_2_17;output CRC_OUT_2_18;output CRC_OUT_2_19;output CRC_OUT_2_2;output CRC_OUT_2_20;output CRC_OUT_2_21;output CRC_OUT_2_22;output CRC_OUT_2_23;output CRC_OUT_2_24;output CRC_OUT_2_25;output CRC_OUT_2_26;output CRC_OUT_2_27;output CRC_OUT_2_28;output CRC_OUT_2_29;output CRC_OUT_2_3;output CRC_OUT_2_30;output CRC_OUT_2_31;output CRC_OUT_2_4;output CRC_OUT_2_5;output CRC_OUT_2_6;output CRC_OUT_2_7;output CRC_OUT_2_8;output CRC_OUT_2_9;output CRC_OUT_3_0;output CRC_OUT_3_1;output CRC_OUT_3_10;output CRC_OUT_3_11;output CRC_OUT_3_12;output CRC_OUT_3_13;output CRC_OUT_3_14;output CRC_OUT_3_15;output CRC_OUT_3_16;output CRC_OUT_3_17;output CRC_OUT_3_18;output CRC_OUT_3_19;output CRC_OUT_3_2;output CRC_OUT_3_20;output CRC_OUT_3_21;output CRC_OUT_3_22;output CRC_OUT_3_23;output CRC_OUT_3_24;output CRC_OUT_3_25;output CRC_OUT_3_26;output CRC_OUT_3_27;output CRC_OUT_3_28;output CRC_OUT_3_29;output CRC_OUT_3_3;output CRC_OUT_3_30;output CRC_OUT_3_31;output CRC_OUT_3_4;output CRC_OUT_3_5;output CRC_OUT_3_6;output CRC_OUT_3_7;output CRC_OUT_3_8;output CRC_OUT_3_9;output CRC_OUT_4_0;output CRC_OUT_4_1;output CRC_OUT_4_10;output CRC_OUT_4_11;output CRC_OUT_4_12;output CRC_OUT_4_13;output CRC_OUT_4_14;output CRC_OUT_4_15;output CRC_OUT_4_16;output CRC_OUT_4_17;output CRC_OUT_4_18;output CRC_OUT_4_19;output CRC_OUT_4_2;output CRC_OUT_4_20;output CRC_OUT_4_21;output CRC_OUT_4_22;output CRC_OUT_4_23;output CRC_OUT_4_24;output CRC_OUT_4_25;output CRC_OUT_4_26;output CRC_OUT_4_27;output CRC_OUT_4_28;output CRC_OUT_4_29;output CRC_OUT_4_3;output CRC_OUT_4_30;output CRC_OUT_4_31;output CRC_OUT_4_4;output CRC_OUT_4_5;output CRC_OUT_4_6;output CRC_OUT_4_7;output CRC_OUT_4_8;output CRC_OUT_4_9;output CRC_OUT_5_0;output CRC_OUT_5_1;output CRC_OUT_5_10;output CRC_OUT_5_11;output CRC_OUT_5_12;output CRC_OUT_5_13;output CRC_OUT_5_14;output CRC_OUT_5_15;output CRC_OUT_5_16;output CRC_OUT_5_17;output CRC_OUT_5_18;output CRC_OUT_5_19;output CRC_OUT_5_2;output CRC_OUT_5_20;output CRC_OUT_5_21;output CRC_OUT_5_22;output CRC_OUT_5_23;output CRC_OUT_5_24;output CRC_OUT_5_25;output CRC_OUT_5_26;output CRC_OUT_5_27;output CRC_OUT_5_28;output CRC_OUT_5_29;output CRC_OUT_5_3;output CRC_OUT_5_30;output CRC_OUT_5_31;output CRC_OUT_5_4;output CRC_OUT_5_5;output CRC_OUT_5_6;output CRC_OUT_5_7;output CRC_OUT_5_8;output CRC_OUT_5_9;output CRC_OUT_6_0;output CRC_OUT_6_1;output CRC_OUT_6_10;output CRC_OUT_6_11;output CRC_OUT_6_12;output CRC_OUT_6_13;output CRC_OUT_6_14;output CRC_OUT_6_15;output CRC_OUT_6_16;output CRC_OUT_6_17;output CRC_OUT_6_18;output CRC_OUT_6_19;output CRC_OUT_6_2;output CRC_OUT_6_20;output CRC_OUT_6_21;output CRC_OUT_6_22;output CRC_OUT_6_23;output CRC_OUT_6_24;output CRC_OUT_6_25;output CRC_OUT_6_26;output CRC_OUT_6_27;output CRC_OUT_6_28;output CRC_OUT_6_29;output CRC_OUT_6_3;output CRC_OUT_6_30;output CRC_OUT_6_31;output CRC_OUT_6_4;output CRC_OUT_6_5;output CRC_OUT_6_6;output CRC_OUT_6_7;output CRC_OUT_6_8;output CRC_OUT_6_9;output CRC_OUT_7_0;output CRC_OUT_7_1;output CRC_OUT_7_10;output CRC_OUT_7_11;output CRC_OUT_7_12;output CRC_OUT_7_13;output CRC_OUT_7_14;output CRC_OUT_7_15;output CRC_OUT_7_16;output CRC_OUT_7_17;output CRC_OUT_7_18;output CRC_OUT_7_19;output CRC_OUT_7_2;output CRC_OUT_7_20;output CRC_OUT_7_21;output CRC_OUT_7_22;output CRC_OUT_7_23;output CRC_OUT_7_24;output CRC_OUT_7_25;output CRC_OUT_7_26;output CRC_OUT_7_27;output CRC_OUT_7_28;output CRC_OUT_7_29;output CRC_OUT_7_3;output CRC_OUT_7_30;output CRC_OUT_7_31;output CRC_OUT_7_4;output CRC_OUT_7_5;output CRC_OUT_7_6;output CRC_OUT_7_7;output CRC_OUT_7_8;output CRC_OUT_7_9;output CRC_OUT_8_0;output CRC_OUT_8_1;output CRC_OUT_8_10;output CRC_OUT_8_11;output CRC_OUT_8_12;output CRC_OUT_8_13;output CRC_OUT_8_14;output CRC_OUT_8_15;output CRC_OUT_8_16;output CRC_OUT_8_17;output CRC_OUT_8_18;output CRC_OUT_8_19;output CRC_OUT_8_2;output CRC_OUT_8_20;output CRC_OUT_8_21;output CRC_OUT_8_22;output CRC_OUT_8_23;output CRC_OUT_8_24;output CRC_OUT_8_25;output CRC_OUT_8_26;output CRC_OUT_8_27;output CRC_OUT_8_28;output CRC_OUT_8_29;output CRC_OUT_8_3;output CRC_OUT_8_30;output CRC_OUT_8_31;output CRC_OUT_8_4;output CRC_OUT_8_5;output CRC_OUT_8_6;output CRC_OUT_8_7;output CRC_OUT_8_8;output CRC_OUT_8_9;output CRC_OUT_9_0;output CRC_OUT_9_1;output CRC_OUT_9_10;output CRC_OUT_9_11;output CRC_OUT_9_12;output CRC_OUT_9_13;output CRC_OUT_9_14;output CRC_OUT_9_15;output CRC_OUT_9_16;output CRC_OUT_9_17;output CRC_OUT_9_18;output CRC_OUT_9_19;output CRC_OUT_9_2;output CRC_OUT_9_20;output CRC_OUT_9_21;output CRC_OUT_9_22;output CRC_OUT_9_23;output CRC_OUT_9_24;output CRC_OUT_9_25;output CRC_OUT_9_26;output CRC_OUT_9_27;output CRC_OUT_9_28;output CRC_OUT_9_29;output CRC_OUT_9_3;output CRC_OUT_9_30;output CRC_OUT_9_31;output CRC_OUT_9_4;output CRC_OUT_9_5;output CRC_OUT_9_6;output CRC_OUT_9_7;output CRC_OUT_9_8;output CRC_OUT_9_9;output DATA_9_0;output DATA_9_1;output DATA_9_10;output DATA_9_11;output DATA_9_12;output DATA_9_13;output DATA_9_14;output DATA_9_15;output DATA_9_16;output DATA_9_17;output DATA_9_18;output DATA_9_19;output DATA_9_2;output DATA_9_20;output DATA_9_21;output DATA_9_22;output DATA_9_23;output DATA_9_24;output DATA_9_25;output DATA_9_26;output DATA_9_27;output DATA_9_28;output DATA_9_29;output DATA_9_3;output DATA_9_30;output DATA_9_31;output DATA_9_4;output DATA_9_5;output DATA_9_6;output DATA_9_7;output DATA_9_8;output DATA_9_9;output test_so;
  wire CRC_OUT_1_31;wire CRC_OUT_1_31_t;wire WX9949;wire WX9949_t;wire WX9947;wire WX9947_t;wire WX9945;wire WX9945_t;wire WX9943;wire WX9943_t;wire WX9941;wire WX9941_t;wire WX9939;wire WX9939_t;wire WX9937;wire WX9937_t;wire WX9935;wire WX9935_t;wire WX9933;wire WX9933_t;wire WX9931;wire WX9931_t;wire WX9929;wire WX9929_t;wire WX9927;wire WX9927_t;wire WX9925;wire WX9925_t;wire WX9923;wire WX9923_t;wire WX9921;wire WX9921_t;wire WX9919;wire WX9919_t;wire WX9917;wire WX9917_t;wire WX9915;wire WX9915_t;wire WX9913;wire WX9913_t;wire WX9911;wire WX9911_t;wire WX9909;wire WX9909_t;wire WX9907;wire WX9907_t;wire WX9905;wire WX9905_t;wire WX9903;wire WX9903_t;wire WX9901;wire WX9901_t;wire WX9899;wire WX9899_t;wire WX9897;wire WX9897_t;wire WX9895;wire WX9895_t;wire WX9893;wire WX9893_t;wire WX9891;wire WX9891_t;wire WX9889;wire WX9889_t;wire WX9887;wire WX9887_t;wire WX9885;wire WX9885_t;wire WX9883;wire WX9883_t;wire WX9881;wire WX9881_t;wire WX9879;wire WX9879_t;wire WX9877;wire WX9877_t;wire WX9875;wire WX9875_t;wire WX9873;wire WX9873_t;wire WX9871;wire WX9871_t;wire WX9869;wire WX9869_t;wire WX9867;wire WX9867_t;wire WX9865;wire WX9865_t;wire WX9863;wire WX9863_t;wire WX9861;wire WX9861_t;wire WX9859;wire WX9859_t;wire WX9857;wire WX9857_t;wire WX9855;wire WX9855_t;wire WX9853;wire WX9853_t;wire WX9851;wire WX9851_t;wire WX9849;wire WX9849_t;wire WX9847;wire WX9847_t;wire WX9845;wire WX9845_t;wire WX9843;wire WX9843_t;wire WX9841;wire WX9841_t;wire WX9839;wire WX9839_t;wire WX9837;wire WX9837_t;wire WX9835;wire WX9835_t;wire WX9833;wire WX9833_t;wire WX9831;wire WX9831_t;wire WX9829;wire WX9829_t;wire WX9827;wire WX9827_t;wire WX9825;wire WX9825_t;wire WX9823;wire WX9823_t;wire WX9821;wire WX9821_t;wire WX9819;wire WX9819_t;wire WX9817;wire WX9817_t;wire WX9815;wire WX9815_t;wire WX9813;wire WX9813_t;wire WX9811;wire WX9811_t;wire WX9809;wire WX9809_t;wire WX9807;wire WX9807_t;wire WX9805;wire WX9805_t;wire WX9803;wire WX9803_t;wire WX9801;wire WX9801_t;wire WX9799;wire WX9799_t;wire WX9797;wire WX9797_t;wire WX9795;wire WX9795_t;wire WX9793;wire WX9793_t;wire WX9791;wire WX9791_t;wire WX9789;wire WX9789_t;wire WX9787;wire WX9787_t;wire WX9785;wire WX9785_t;wire WX9783;wire WX9783_t;wire WX9781;wire WX9781_t;wire WX9779;wire WX9779_t;wire WX9777;wire WX9777_t;wire WX9775;wire WX9775_t;wire WX9773;wire WX9773_t;wire WX9771;wire WX9771_t;wire WX9769;wire WX9769_t;wire WX9767;wire WX9767_t;wire WX9765;wire WX9765_t;wire WX9763;wire WX9763_t;wire WX9761;wire WX9761_t;wire WX9759;wire WX9759_t;wire WX9757;wire WX9757_t;wire WX9755;wire WX9755_t;wire WX9753;wire WX9753_t;wire WX9751;wire WX9751_t;wire WX9749;wire WX9749_t;wire WX9747;wire WX9747_t;wire WX9745;wire WX9745_t;wire WX9743;wire WX9743_t;wire WX9741;wire WX9741_t;wire WX9739;wire WX9739_t;wire WX9737;wire WX9737_t;wire WX9735;wire WX9735_t;wire WX9733;wire WX9733_t;wire WX9731;wire WX9731_t;wire WX9729;wire WX9729_t;wire WX9727;wire WX9727_t;wire WX9725;wire WX9725_t;wire WX9723;wire WX9723_t;wire WX9721;wire WX9721_t;wire WX9719;wire WX9719_t;wire WX9717;wire WX9717_t;wire WX9715;wire WX9715_t;wire WX9713;wire WX9713_t;wire WX9711;wire WX9711_t;wire WX9709;wire WX9709_t;wire WX9707;wire WX9707_t;wire WX9705;wire WX9705_t;wire WX9703;wire WX9703_t;wire WX9701;wire WX9701_t;wire WX9699;wire WX9699_t;wire WX9697;wire WX9697_t;wire WX9695;wire WX9695_t;wire WX9597;wire WX9597_t;wire WX9595;wire WX9595_t;wire WX9593;wire WX9593_t;wire WX9591;wire WX9591_t;wire WX9589;wire WX9589_t;wire WX9587;wire WX9587_t;wire WX9585;wire WX9585_t;wire WX9583;wire WX9583_t;wire WX9581;wire WX9581_t;wire WX9579;wire WX9579_t;wire WX9577;wire WX9577_t;wire WX9575;wire WX9575_t;wire WX9573;wire WX9573_t;wire WX9571;wire WX9571_t;wire WX9569;wire WX9569_t;wire WX9567;wire WX9567_t;wire WX9565;wire WX9565_t;wire WX9563;wire WX9563_t;wire WX9561;wire WX9561_t;wire WX9559;wire WX9559_t;wire WX9557;wire WX9557_t;wire WX9555;wire WX9555_t;wire WX9553;wire WX9553_t;wire WX9551;wire WX9551_t;wire WX9549;wire WX9549_t;wire WX9547;wire WX9547_t;wire WX9545;wire WX9545_t;wire WX9543;wire WX9543_t;wire WX9541;wire WX9541_t;wire WX9539;wire WX9539_t;wire WX9537;wire WX9537_t;wire WX9535;wire WX9535_t;wire WX9084;wire WX9084_t;wire WX9082;wire WX9082_t;wire WX9080;wire WX9080_t;wire WX9078;wire WX9078_t;wire WX9076;wire WX9076_t;wire WX9074;wire WX9074_t;wire WX9072;wire WX9072_t;wire WX9070;wire WX9070_t;wire WX9068;wire WX9068_t;wire WX9066;wire WX9066_t;wire WX9064;wire WX9064_t;wire WX9062;wire WX9062_t;wire WX9060;wire WX9060_t;wire WX9058;wire WX9058_t;wire WX9056;wire WX9056_t;wire WX9054;wire WX9054_t;wire WX9052;wire WX9052_t;wire WX9050;wire WX9050_t;wire WX9048;wire WX9048_t;wire WX9046;wire WX9046_t;wire WX9044;wire WX9044_t;wire WX9042;wire WX9042_t;wire WX9040;wire WX9040_t;wire WX9038;wire WX9038_t;wire WX9036;wire WX9036_t;wire WX9034;wire WX9034_t;wire WX9032;wire WX9032_t;wire WX9030;wire WX9030_t;wire WX9028;wire WX9028_t;wire WX9026;wire WX9026_t;wire WX9024;wire WX9024_t;wire WX9022;wire WX9022_t;wire WX898;wire WX898_t;wire WX896;wire WX896_t;wire WX894;wire WX894_t;wire WX892;wire WX892_t;wire WX890;wire WX890_t;wire WX888;wire WX888_t;wire WX886;wire WX886_t;wire WX884;wire WX884_t;wire WX882;wire WX882_t;wire WX880;wire WX880_t;wire WX878;wire WX878_t;wire WX876;wire WX876_t;wire WX874;wire WX874_t;wire WX872;wire WX872_t;wire WX870;wire WX870_t;wire WX868;wire WX868_t;wire WX866;wire WX866_t;wire WX8656;wire WX8656_t;wire WX8654;wire WX8654_t;wire WX8652;wire WX8652_t;wire WX8650;wire WX8650_t;wire WX8648;wire WX8648_t;wire WX8646;wire WX8646_t;wire WX8644;wire WX8644_t;wire WX8642;wire WX8642_t;wire WX8640;wire WX8640_t;wire WX864;wire WX864_t;wire WX8638;wire WX8638_t;wire WX8636;wire WX8636_t;wire WX8634;wire WX8634_t;wire WX8632;wire WX8632_t;wire WX8630;wire WX8630_t;wire WX8628;wire WX8628_t;wire WX8626;wire WX8626_t;wire WX8624;wire WX8624_t;wire WX8622;wire WX8622_t;wire WX8620;wire WX8620_t;wire WX862;wire WX862_t;wire WX8618;wire WX8618_t;wire WX8616;wire WX8616_t;wire WX8614;wire WX8614_t;wire WX8612;wire WX8612_t;wire WX8610;wire WX8610_t;wire WX8608;wire WX8608_t;wire WX8606;wire WX8606_t;wire WX8604;wire WX8604_t;wire WX8602;wire WX8602_t;wire WX8600;wire WX8600_t;wire WX860;wire WX860_t;wire WX8598;wire WX8598_t;wire WX8596;wire WX8596_t;wire WX8594;wire WX8594_t;wire WX8592;wire WX8592_t;wire WX8590;wire WX8590_t;wire WX8588;wire WX8588_t;wire WX8586;wire WX8586_t;wire WX8584;wire WX8584_t;wire WX8582;wire WX8582_t;wire WX8580;wire WX8580_t;wire WX858;wire WX858_t;wire WX8578;wire WX8578_t;wire WX8576;wire WX8576_t;wire WX8574;wire WX8574_t;wire WX8572;wire WX8572_t;wire WX8570;wire WX8570_t;wire WX8568;wire WX8568_t;wire WX8566;wire WX8566_t;wire WX8564;wire WX8564_t;wire WX8562;wire WX8562_t;wire WX8560;wire WX8560_t;wire WX856;wire WX856_t;wire WX8558;wire WX8558_t;wire WX8556;wire WX8556_t;wire WX8554;wire WX8554_t;wire WX8552;wire WX8552_t;wire WX8550;wire WX8550_t;wire WX8548;wire WX8548_t;wire WX8546;wire WX8546_t;wire WX8544;wire WX8544_t;wire WX8542;wire WX8542_t;wire WX8540;wire WX8540_t;wire WX854;wire WX854_t;wire WX8538;wire WX8538_t;wire WX8536;wire WX8536_t;wire WX8534;wire WX8534_t;wire WX8532;wire WX8532_t;wire WX8530;wire WX8530_t;wire WX8528;wire WX8528_t;wire WX8526;wire WX8526_t;wire WX8524;wire WX8524_t;wire WX8522;wire WX8522_t;wire WX8520;wire WX8520_t;wire WX852;wire WX852_t;wire WX8518;wire WX8518_t;wire WX8516;wire WX8516_t;wire WX8514;wire WX8514_t;wire WX8512;wire WX8512_t;wire WX8510;wire WX8510_t;wire WX8508;wire WX8508_t;wire WX8506;wire WX8506_t;wire WX8504;wire WX8504_t;wire WX8502;wire WX8502_t;wire WX8500;wire WX8500_t;wire WX850;wire WX850_t;wire WX8498;wire WX8498_t;wire WX8496;wire WX8496_t;wire WX8494;wire WX8494_t;wire WX8492;wire WX8492_t;wire WX8490;wire WX8490_t;wire WX8488;wire WX8488_t;wire WX8486;wire WX8486_t;wire WX8484;wire WX8484_t;wire WX8482;wire WX8482_t;wire WX8480;wire WX8480_t;wire WX848;wire WX848_t;wire WX8478;wire WX8478_t;wire WX8476;wire WX8476_t;wire WX8474;wire WX8474_t;wire WX8472;wire WX8472_t;wire WX8470;wire WX8470_t;wire WX8468;wire WX8468_t;wire WX8466;wire WX8466_t;wire WX8464;wire WX8464_t;wire n3205;wire n3205_t;wire WX8462;wire WX8462_t;wire n3206;wire n3206_t;wire WX8460;wire WX8460_t;wire n3207;wire n3207_t;wire WX846;wire WX846_t;wire WX8458;wire WX8458_t;wire n3208;wire n3208_t;wire WX8456;wire WX8456_t;wire n3209;wire n3209_t;wire WX8454;wire WX8454_t;wire n3210;wire n3210_t;wire WX8452;wire WX8452_t;wire n3211;wire n3211_t;wire WX8450;wire WX8450_t;wire n3212;wire n3212_t;wire WX8448;wire WX8448_t;wire n3213;wire n3213_t;wire WX8446;wire WX8446_t;wire n3214;wire n3214_t;wire WX8444;wire WX8444_t;wire n3215;wire n3215_t;wire WX8442;wire WX8442_t;wire n3216;wire n3216_t;wire WX8440;wire WX8440_t;wire n3217;wire n3217_t;wire WX844;wire WX844_t;wire WX8438;wire WX8438_t;wire n3218;wire n3218_t;wire WX8436;wire WX8436_t;wire n3219;wire n3219_t;wire WX8434;wire WX8434_t;wire n3220;wire n3220_t;wire WX8432;wire WX8432_t;wire WX8430;wire WX8430_t;wire WX8428;wire WX8428_t;wire WX8426;wire WX8426_t;wire WX8424;wire WX8424_t;wire WX8422;wire WX8422_t;wire WX8420;wire WX8420_t;wire WX842;wire WX842_t;wire WX8418;wire WX8418_t;wire WX8416;wire WX8416_t;wire WX8414;wire WX8414_t;wire WX8412;wire WX8412_t;wire WX8410;wire WX8410_t;wire WX8408;wire WX8408_t;wire WX8406;wire WX8406_t;wire WX8404;wire WX8404_t;wire WX8402;wire WX8402_t;wire WX840;wire WX840_t;wire WX838;wire WX838_t;wire WX836;wire WX836_t;wire WX834;wire WX834_t;wire WX832;wire WX832_t;wire WX8304;wire WX8304_t;wire WX8302;wire WX8302_t;wire WX8300;wire WX8300_t;wire WX830;wire WX830_t;wire WX8298;wire WX8298_t;wire WX8296;wire WX8296_t;wire WX8294;wire WX8294_t;wire WX8292;wire WX8292_t;wire WX8290;wire WX8290_t;wire WX8288;wire WX8288_t;wire WX8286;wire WX8286_t;wire WX8284;wire WX8284_t;wire WX8282;wire WX8282_t;wire WX8280;wire WX8280_t;wire WX828;wire WX828_t;wire WX8278;wire WX8278_t;wire WX8276;wire WX8276_t;wire WX8274;wire WX8274_t;wire WX8272;wire WX8272_t;wire WX8270;wire WX8270_t;wire WX8268;wire WX8268_t;wire WX8266;wire WX8266_t;wire WX8264;wire WX8264_t;wire WX8262;wire WX8262_t;wire WX8260;wire WX8260_t;wire WX826;wire WX826_t;wire WX8258;wire WX8258_t;wire WX8256;wire WX8256_t;wire WX8254;wire WX8254_t;wire WX8252;wire WX8252_t;wire WX8250;wire WX8250_t;wire WX8248;wire WX8248_t;wire WX8246;wire WX8246_t;wire WX8244;wire WX8244_t;wire WX8242;wire WX8242_t;wire WX824;wire WX824_t;wire WX822;wire WX822_t;wire WX820;wire WX820_t;wire WX818;wire WX818_t;wire WX816;wire WX816_t;wire WX814;wire WX814_t;wire WX812;wire WX812_t;wire WX810;wire WX810_t;wire WX808;wire WX808_t;wire WX806;wire WX806_t;wire WX804;wire WX804_t;wire WX802;wire WX802_t;wire WX800;wire WX800_t;wire WX798;wire WX798_t;wire WX796;wire WX796_t;wire WX794;wire WX794_t;wire WX792;wire WX792_t;wire WX790;wire WX790_t;wire WX788;wire WX788_t;wire WX786;wire WX786_t;wire WX784;wire WX784_t;wire WX782;wire WX782_t;wire WX780;wire WX780_t;wire WX7791;wire WX7791_t;wire WX7789;wire WX7789_t;wire WX7787;wire WX7787_t;wire WX7785;wire WX7785_t;wire WX7783;wire WX7783_t;wire WX7781;wire WX7781_t;wire WX778;wire WX778_t;wire WX7779;wire WX7779_t;wire WX7777;wire WX7777_t;wire WX7775;wire WX7775_t;wire WX7773;wire WX7773_t;wire WX7771;wire WX7771_t;wire WX7769;wire WX7769_t;wire WX7767;wire WX7767_t;wire WX7765;wire WX7765_t;wire WX7763;wire WX7763_t;wire WX7761;wire WX7761_t;wire WX776;wire WX776_t;wire WX7759;wire WX7759_t;wire WX7757;wire WX7757_t;wire WX7755;wire WX7755_t;wire WX7753;wire WX7753_t;wire WX7751;wire WX7751_t;wire WX7749;wire WX7749_t;wire WX7747;wire WX7747_t;wire WX7745;wire WX7745_t;wire WX7743;wire WX7743_t;wire WX7741;wire WX7741_t;wire WX774;wire WX774_t;wire WX7739;wire WX7739_t;wire WX7737;wire WX7737_t;wire WX7735;wire WX7735_t;wire WX7733;wire WX7733_t;wire WX7731;wire WX7731_t;wire WX7729;wire WX7729_t;wire WX772;wire WX772_t;wire WX770;wire WX770_t;wire WX768;wire WX768_t;wire WX766;wire WX766_t;wire WX764;wire WX764_t;wire WX762;wire WX762_t;wire WX760;wire WX760_t;wire WX758;wire WX758_t;wire WX756;wire WX756_t;wire WX754;wire WX754_t;wire WX752;wire WX752_t;wire WX750;wire WX750_t;wire WX748;wire WX748_t;wire WX746;wire WX746_t;wire WX744;wire WX744_t;wire WX742;wire WX742_t;wire WX740;wire WX740_t;wire WX738;wire WX738_t;wire WX7363;wire WX7363_t;wire WX7361;wire WX7361_t;wire WX736;wire WX736_t;wire WX7359;wire WX7359_t;wire WX7357;wire WX7357_t;wire WX7355;wire WX7355_t;wire WX7353;wire WX7353_t;wire WX7351;wire WX7351_t;wire WX7349;wire WX7349_t;wire WX7347;wire WX7347_t;wire WX7345;wire WX7345_t;wire WX7343;wire WX7343_t;wire WX7341;wire WX7341_t;wire WX734;wire WX734_t;wire WX7339;wire WX7339_t;wire WX7337;wire WX7337_t;wire WX7335;wire WX7335_t;wire WX7333;wire WX7333_t;wire WX7331;wire WX7331_t;wire WX7329;wire WX7329_t;wire WX7327;wire WX7327_t;wire WX7325;wire WX7325_t;wire WX7323;wire WX7323_t;wire WX7321;wire WX7321_t;wire WX732;wire WX732_t;wire WX7319;wire WX7319_t;wire WX7317;wire WX7317_t;wire WX7315;wire WX7315_t;wire WX7313;wire WX7313_t;wire WX7311;wire WX7311_t;wire WX7309;wire WX7309_t;wire WX7307;wire WX7307_t;wire WX7305;wire WX7305_t;wire WX7303;wire WX7303_t;wire WX7301;wire WX7301_t;wire WX730;wire WX730_t;wire WX7299;wire WX7299_t;wire WX7297;wire WX7297_t;wire WX7295;wire WX7295_t;wire WX7293;wire WX7293_t;wire WX7291;wire WX7291_t;wire WX7289;wire WX7289_t;wire WX7287;wire WX7287_t;wire WX7285;wire WX7285_t;wire WX7283;wire WX7283_t;wire WX7281;wire WX7281_t;wire WX728;wire WX728_t;wire WX7279;wire WX7279_t;wire WX7277;wire WX7277_t;wire WX7275;wire WX7275_t;wire WX7273;wire WX7273_t;wire WX7271;wire WX7271_t;wire WX7269;wire WX7269_t;wire WX7267;wire WX7267_t;wire WX7265;wire WX7265_t;wire WX7263;wire WX7263_t;wire WX7261;wire WX7261_t;wire WX726;wire WX726_t;wire WX7259;wire WX7259_t;wire WX7257;wire WX7257_t;wire WX7255;wire WX7255_t;wire WX7253;wire WX7253_t;wire WX7251;wire WX7251_t;wire WX7249;wire WX7249_t;wire WX7247;wire WX7247_t;wire WX7245;wire WX7245_t;wire WX7243;wire WX7243_t;wire WX7241;wire WX7241_t;wire WX724;wire WX724_t;wire WX7239;wire WX7239_t;wire WX7237;wire WX7237_t;wire WX7235;wire WX7235_t;wire WX7233;wire WX7233_t;wire WX7231;wire WX7231_t;wire WX7229;wire WX7229_t;wire WX7227;wire WX7227_t;wire WX7225;wire WX7225_t;wire WX7223;wire WX7223_t;wire WX7221;wire WX7221_t;wire WX722;wire WX722_t;wire WX7219;wire WX7219_t;wire WX7217;wire WX7217_t;wire WX7215;wire WX7215_t;wire WX7213;wire WX7213_t;wire WX7211;wire WX7211_t;wire WX7209;wire WX7209_t;wire WX7207;wire WX7207_t;wire WX7205;wire WX7205_t;wire WX7203;wire WX7203_t;wire WX7201;wire WX7201_t;wire WX720;wire WX720_t;wire WX7199;wire WX7199_t;wire WX7197;wire WX7197_t;wire WX7195;wire WX7195_t;wire WX7193;wire WX7193_t;wire WX7191;wire WX7191_t;wire WX7189;wire WX7189_t;wire WX7187;wire WX7187_t;wire WX7185;wire WX7185_t;wire WX7183;wire WX7183_t;wire WX7181;wire WX7181_t;wire WX718;wire WX718_t;wire WX7179;wire WX7179_t;wire WX7177;wire WX7177_t;wire WX7175;wire WX7175_t;wire WX7173;wire WX7173_t;wire WX7171;wire WX7171_t;wire n3221;wire n3221_t;wire WX7169;wire WX7169_t;wire n3222;wire n3222_t;wire WX7167;wire WX7167_t;wire n3223;wire n3223_t;wire WX7165;wire WX7165_t;wire n3224;wire n3224_t;wire WX7163;wire WX7163_t;wire n3225;wire n3225_t;wire WX7161;wire WX7161_t;wire n3226;wire n3226_t;wire WX716;wire WX716_t;wire WX7159;wire WX7159_t;wire n3227;wire n3227_t;wire WX7157;wire WX7157_t;wire n3228;wire n3228_t;wire WX7155;wire WX7155_t;wire n3229;wire n3229_t;wire WX7153;wire WX7153_t;wire n3230;wire n3230_t;wire WX7151;wire WX7151_t;wire n3231;wire n3231_t;wire WX7149;wire WX7149_t;wire n3232;wire n3232_t;wire WX7147;wire WX7147_t;wire n3233;wire n3233_t;wire WX7145;wire WX7145_t;wire n3234;wire n3234_t;wire WX7143;wire WX7143_t;wire n3235;wire n3235_t;wire WX7141;wire WX7141_t;wire n3236;wire n3236_t;wire WX714;wire WX714_t;wire WX7139;wire WX7139_t;wire WX7137;wire WX7137_t;wire WX7135;wire WX7135_t;wire WX7133;wire WX7133_t;wire WX7131;wire WX7131_t;wire WX7129;wire WX7129_t;wire WX7127;wire WX7127_t;wire WX7125;wire WX7125_t;wire WX7123;wire WX7123_t;wire WX7121;wire WX7121_t;wire WX712;wire WX712_t;wire WX7119;wire WX7119_t;wire WX7117;wire WX7117_t;wire WX7115;wire WX7115_t;wire WX7113;wire WX7113_t;wire WX7111;wire WX7111_t;wire WX7109;wire WX7109_t;wire WX710;wire WX710_t;wire WX708;wire WX708_t;wire WX706;wire WX706_t;wire WX704;wire WX704_t;wire WX702;wire WX702_t;wire WX7011;wire WX7011_t;wire WX7009;wire WX7009_t;wire WX7007;wire WX7007_t;wire WX7005;wire WX7005_t;wire WX7003;wire WX7003_t;wire WX7001;wire WX7001_t;wire WX700;wire WX700_t;wire WX6999;wire WX6999_t;wire WX6997;wire WX6997_t;wire WX6995;wire WX6995_t;wire WX6993;wire WX6993_t;wire WX6991;wire WX6991_t;wire WX6989;wire WX6989_t;wire WX6987;wire WX6987_t;wire WX6985;wire WX6985_t;wire WX6983;wire WX6983_t;wire WX6981;wire WX6981_t;wire WX698;wire WX698_t;wire WX6979;wire WX6979_t;wire WX6977;wire WX6977_t;wire WX6975;wire WX6975_t;wire WX6973;wire WX6973_t;wire WX6971;wire WX6971_t;wire WX6969;wire WX6969_t;wire WX6967;wire WX6967_t;wire WX6965;wire WX6965_t;wire WX6963;wire WX6963_t;wire WX6961;wire WX6961_t;wire WX696;wire WX696_t;wire WX6959;wire WX6959_t;wire WX6957;wire WX6957_t;wire WX6955;wire WX6955_t;wire WX6953;wire WX6953_t;wire WX6951;wire WX6951_t;wire WX6949;wire WX6949_t;wire WX694;wire WX694_t;wire WX692;wire WX692_t;wire WX690;wire WX690_t;wire WX688;wire WX688_t;wire WX686;wire WX686_t;wire WX684;wire WX684_t;wire WX682;wire WX682_t;wire WX680;wire WX680_t;wire WX678;wire WX678_t;wire WX676;wire WX676_t;wire WX674;wire WX674_t;wire WX672;wire WX672_t;wire WX670;wire WX670_t;wire WX668;wire WX668_t;wire WX666;wire WX666_t;wire WX664;wire WX664_t;wire WX662;wire WX662_t;wire WX660;wire WX660_t;wire WX658;wire WX658_t;wire WX656;wire WX656_t;wire WX654;wire WX654_t;wire WX652;wire WX652_t;wire WX650;wire WX650_t;wire WX6498;wire WX6498_t;wire WX6496;wire WX6496_t;wire WX6494;wire WX6494_t;wire WX6492;wire WX6492_t;wire WX6490;wire WX6490_t;wire WX6488;wire WX6488_t;wire WX6486;wire WX6486_t;wire WX6484;wire WX6484_t;wire WX6482;wire WX6482_t;wire WX6480;wire WX6480_t;wire WX648;wire WX648_t;wire WX6478;wire WX6478_t;wire WX6476;wire WX6476_t;wire WX6474;wire WX6474_t;wire WX6472;wire WX6472_t;wire WX6470;wire WX6470_t;wire WX6468;wire WX6468_t;wire WX6466;wire WX6466_t;wire WX6464;wire WX6464_t;wire WX6462;wire WX6462_t;wire WX6460;wire WX6460_t;wire WX646;wire WX646_t;wire WX6458;wire WX6458_t;wire WX6456;wire WX6456_t;wire WX6454;wire WX6454_t;wire WX6452;wire WX6452_t;wire WX6450;wire WX6450_t;wire WX6448;wire WX6448_t;wire WX6446;wire WX6446_t;wire WX6444;wire WX6444_t;wire WX6442;wire WX6442_t;wire WX6440;wire WX6440_t;wire WX644;wire WX644_t;wire WX6438;wire WX6438_t;wire WX6436;wire WX6436_t;wire WX6070;wire WX6070_t;wire WX6068;wire WX6068_t;wire WX6066;wire WX6066_t;wire WX6064;wire WX6064_t;wire WX6062;wire WX6062_t;wire WX6060;wire WX6060_t;wire WX6058;wire WX6058_t;wire WX6056;wire WX6056_t;wire WX6054;wire WX6054_t;wire WX6052;wire WX6052_t;wire WX6050;wire WX6050_t;wire WX6048;wire WX6048_t;wire WX6046;wire WX6046_t;wire WX6044;wire WX6044_t;wire WX6042;wire WX6042_t;wire WX6040;wire WX6040_t;wire WX6038;wire WX6038_t;wire WX6036;wire WX6036_t;wire WX6034;wire WX6034_t;wire WX6032;wire WX6032_t;wire WX6030;wire WX6030_t;wire WX6028;wire WX6028_t;wire WX6026;wire WX6026_t;wire WX6024;wire WX6024_t;wire WX6022;wire WX6022_t;wire WX6020;wire WX6020_t;wire WX6018;wire WX6018_t;wire WX6016;wire WX6016_t;wire WX6014;wire WX6014_t;wire WX6012;wire WX6012_t;wire WX6010;wire WX6010_t;wire WX6008;wire WX6008_t;wire WX6006;wire WX6006_t;wire WX6004;wire WX6004_t;wire WX6002;wire WX6002_t;wire WX6000;wire WX6000_t;wire WX5998;wire WX5998_t;wire WX5996;wire WX5996_t;wire WX5994;wire WX5994_t;wire WX5992;wire WX5992_t;wire WX5990;wire WX5990_t;wire WX5988;wire WX5988_t;wire WX5986;wire WX5986_t;wire WX5984;wire WX5984_t;wire WX5982;wire WX5982_t;wire WX5980;wire WX5980_t;wire WX5978;wire WX5978_t;wire WX5976;wire WX5976_t;wire WX5974;wire WX5974_t;wire WX5972;wire WX5972_t;wire WX5970;wire WX5970_t;wire WX5968;wire WX5968_t;wire WX5966;wire WX5966_t;wire WX5964;wire WX5964_t;wire WX5962;wire WX5962_t;wire WX5960;wire WX5960_t;wire WX5958;wire WX5958_t;wire WX5956;wire WX5956_t;wire WX5954;wire WX5954_t;wire WX5952;wire WX5952_t;wire WX5950;wire WX5950_t;wire WX5948;wire WX5948_t;wire WX5946;wire WX5946_t;wire WX5944;wire WX5944_t;wire WX5942;wire WX5942_t;wire WX5940;wire WX5940_t;wire WX5938;wire WX5938_t;wire WX5936;wire WX5936_t;wire WX5934;wire WX5934_t;wire WX5932;wire WX5932_t;wire WX5930;wire WX5930_t;wire WX5928;wire WX5928_t;wire WX5926;wire WX5926_t;wire WX5924;wire WX5924_t;wire WX5922;wire WX5922_t;wire WX5920;wire WX5920_t;wire WX5918;wire WX5918_t;wire WX5916;wire WX5916_t;wire WX5914;wire WX5914_t;wire WX5912;wire WX5912_t;wire WX5910;wire WX5910_t;wire WX5908;wire WX5908_t;wire WX5906;wire WX5906_t;wire WX5904;wire WX5904_t;wire WX5902;wire WX5902_t;wire WX5900;wire WX5900_t;wire WX5898;wire WX5898_t;wire WX5896;wire WX5896_t;wire WX5894;wire WX5894_t;wire WX5892;wire WX5892_t;wire WX5890;wire WX5890_t;wire WX5888;wire WX5888_t;wire WX5886;wire WX5886_t;wire WX5884;wire WX5884_t;wire WX5882;wire WX5882_t;wire WX5880;wire WX5880_t;wire WX5878;wire WX5878_t;wire n3237;wire n3237_t;wire WX5876;wire WX5876_t;wire n3238;wire n3238_t;wire WX5874;wire WX5874_t;wire n3239;wire n3239_t;wire WX5872;wire WX5872_t;wire n3240;wire n3240_t;wire WX5870;wire WX5870_t;wire n3241;wire n3241_t;wire WX5868;wire WX5868_t;wire n3242;wire n3242_t;wire WX5866;wire WX5866_t;wire n3243;wire n3243_t;wire WX5864;wire WX5864_t;wire n3244;wire n3244_t;wire WX5862;wire WX5862_t;wire n3245;wire n3245_t;wire WX5860;wire WX5860_t;wire n3246;wire n3246_t;wire WX5858;wire WX5858_t;wire n3247;wire n3247_t;wire WX5856;wire WX5856_t;wire n3248;wire n3248_t;wire WX5854;wire WX5854_t;wire n3249;wire n3249_t;wire WX5852;wire WX5852_t;wire n3250;wire n3250_t;wire WX5850;wire WX5850_t;wire n3251;wire n3251_t;wire WX5848;wire WX5848_t;wire n3252;wire n3252_t;wire WX5846;wire WX5846_t;wire WX5844;wire WX5844_t;wire WX5842;wire WX5842_t;wire WX5840;wire WX5840_t;wire WX5838;wire WX5838_t;wire WX5836;wire WX5836_t;wire WX5834;wire WX5834_t;wire WX5832;wire WX5832_t;wire WX5830;wire WX5830_t;wire WX5828;wire WX5828_t;wire WX5826;wire WX5826_t;wire WX5824;wire WX5824_t;wire WX5822;wire WX5822_t;wire WX5820;wire WX5820_t;wire WX5818;wire WX5818_t;wire WX5816;wire WX5816_t;wire WX5718;wire WX5718_t;wire WX5716;wire WX5716_t;wire WX5714;wire WX5714_t;wire WX5712;wire WX5712_t;wire WX5710;wire WX5710_t;wire WX5708;wire WX5708_t;wire WX5706;wire WX5706_t;wire WX5704;wire WX5704_t;wire WX5702;wire WX5702_t;wire WX5700;wire WX5700_t;wire WX5698;wire WX5698_t;wire WX5696;wire WX5696_t;wire WX5694;wire WX5694_t;wire WX5692;wire WX5692_t;wire WX5690;wire WX5690_t;wire WX5688;wire WX5688_t;wire WX5686;wire WX5686_t;wire WX5684;wire WX5684_t;wire WX5682;wire WX5682_t;wire WX5680;wire WX5680_t;wire WX5678;wire WX5678_t;wire WX5676;wire WX5676_t;wire WX5674;wire WX5674_t;wire WX5672;wire WX5672_t;wire WX5670;wire WX5670_t;wire WX5668;wire WX5668_t;wire WX5666;wire WX5666_t;wire WX5664;wire WX5664_t;wire WX5662;wire WX5662_t;wire WX5660;wire WX5660_t;wire WX5658;wire WX5658_t;wire WX5656;wire WX5656_t;wire WX546;wire WX546_t;wire WX544;wire WX544_t;wire WX542;wire WX542_t;wire WX540;wire WX540_t;wire WX538;wire WX538_t;wire WX536;wire WX536_t;wire WX534;wire WX534_t;wire WX532;wire WX532_t;wire WX530;wire WX530_t;wire WX528;wire WX528_t;wire WX526;wire WX526_t;wire WX524;wire WX524_t;wire WX522;wire WX522_t;wire WX5205;wire WX5205_t;wire WX5203;wire WX5203_t;wire WX5201;wire WX5201_t;wire WX520;wire WX520_t;wire WX5199;wire WX5199_t;wire WX5197;wire WX5197_t;wire WX5195;wire WX5195_t;wire WX5193;wire WX5193_t;wire WX5191;wire WX5191_t;wire WX5189;wire WX5189_t;wire WX5187;wire WX5187_t;wire WX5185;wire WX5185_t;wire WX5183;wire WX5183_t;wire WX5181;wire WX5181_t;wire WX518;wire WX518_t;wire WX5179;wire WX5179_t;wire WX5177;wire WX5177_t;wire WX5175;wire WX5175_t;wire WX5173;wire WX5173_t;wire WX5171;wire WX5171_t;wire WX5169;wire WX5169_t;wire WX5167;wire WX5167_t;wire WX5165;wire WX5165_t;wire WX5163;wire WX5163_t;wire WX5161;wire WX5161_t;wire WX516;wire WX516_t;wire WX5159;wire WX5159_t;wire WX5157;wire WX5157_t;wire WX5155;wire WX5155_t;wire WX5153;wire WX5153_t;wire WX5151;wire WX5151_t;wire WX5149;wire WX5149_t;wire WX5147;wire WX5147_t;wire WX5145;wire WX5145_t;wire WX5143;wire WX5143_t;wire WX514;wire WX514_t;wire WX512;wire WX512_t;wire WX510;wire WX510_t;wire WX508;wire WX508_t;wire WX506;wire WX506_t;wire WX504;wire WX504_t;wire WX502;wire WX502_t;wire WX500;wire WX500_t;wire WX498;wire WX498_t;wire WX496;wire WX496_t;wire WX494;wire WX494_t;wire WX492;wire WX492_t;wire WX490;wire WX490_t;wire WX488;wire WX488_t;wire WX486;wire WX486_t;wire WX484;wire WX484_t;wire WX4777;wire WX4777_t;wire WX4775;wire WX4775_t;wire WX4773;wire WX4773_t;wire WX4771;wire WX4771_t;wire WX4769;wire WX4769_t;wire WX4767;wire WX4767_t;wire WX4765;wire WX4765_t;wire WX4763;wire WX4763_t;wire WX4761;wire WX4761_t;wire WX4759;wire WX4759_t;wire WX4757;wire WX4757_t;wire WX4755;wire WX4755_t;wire WX4753;wire WX4753_t;wire WX4751;wire WX4751_t;wire WX4749;wire WX4749_t;wire WX4747;wire WX4747_t;wire WX4745;wire WX4745_t;wire WX4743;wire WX4743_t;wire WX4741;wire WX4741_t;wire WX4739;wire WX4739_t;wire WX4737;wire WX4737_t;wire WX4735;wire WX4735_t;wire WX4733;wire WX4733_t;wire WX4731;wire WX4731_t;wire WX4729;wire WX4729_t;wire WX4727;wire WX4727_t;wire WX4725;wire WX4725_t;wire WX4723;wire WX4723_t;wire WX4721;wire WX4721_t;wire WX4719;wire WX4719_t;wire WX4717;wire WX4717_t;wire WX4715;wire WX4715_t;wire WX4713;wire WX4713_t;wire WX4711;wire WX4711_t;wire WX4709;wire WX4709_t;wire WX4707;wire WX4707_t;wire WX4705;wire WX4705_t;wire WX4703;wire WX4703_t;wire WX4701;wire WX4701_t;wire WX4699;wire WX4699_t;wire WX4697;wire WX4697_t;wire WX4695;wire WX4695_t;wire WX4693;wire WX4693_t;wire WX4691;wire WX4691_t;wire WX4689;wire WX4689_t;wire WX4687;wire WX4687_t;wire WX4685;wire WX4685_t;wire WX4683;wire WX4683_t;wire WX4681;wire WX4681_t;wire WX4679;wire WX4679_t;wire WX4677;wire WX4677_t;wire WX4675;wire WX4675_t;wire WX4673;wire WX4673_t;wire WX4671;wire WX4671_t;wire WX4669;wire WX4669_t;wire WX4667;wire WX4667_t;wire WX4665;wire WX4665_t;wire WX4663;wire WX4663_t;wire WX4661;wire WX4661_t;wire WX4659;wire WX4659_t;wire WX4657;wire WX4657_t;wire WX4655;wire WX4655_t;wire WX4653;wire WX4653_t;wire WX4651;wire WX4651_t;wire WX4649;wire WX4649_t;wire WX4647;wire WX4647_t;wire WX4645;wire WX4645_t;wire WX4643;wire WX4643_t;wire WX4641;wire WX4641_t;wire WX4639;wire WX4639_t;wire WX4637;wire WX4637_t;wire WX4635;wire WX4635_t;wire WX4633;wire WX4633_t;wire WX4631;wire WX4631_t;wire WX4629;wire WX4629_t;wire WX4627;wire WX4627_t;wire WX4625;wire WX4625_t;wire WX4623;wire WX4623_t;wire WX4621;wire WX4621_t;wire WX4619;wire WX4619_t;wire WX4617;wire WX4617_t;wire WX4615;wire WX4615_t;wire WX4613;wire WX4613_t;wire WX4611;wire WX4611_t;wire WX4609;wire WX4609_t;wire WX4607;wire WX4607_t;wire WX4605;wire WX4605_t;wire WX4603;wire WX4603_t;wire WX4601;wire WX4601_t;wire WX4599;wire WX4599_t;wire WX4597;wire WX4597_t;wire WX4595;wire WX4595_t;wire WX4593;wire WX4593_t;wire WX4591;wire WX4591_t;wire WX4589;wire WX4589_t;wire WX4587;wire WX4587_t;wire WX4585;wire WX4585_t;wire n3253;wire n3253_t;wire WX4583;wire WX4583_t;wire n3254;wire n3254_t;wire WX4581;wire WX4581_t;wire n3255;wire n3255_t;wire WX4579;wire WX4579_t;wire n3256;wire n3256_t;wire WX4577;wire WX4577_t;wire n3257;wire n3257_t;wire WX4575;wire WX4575_t;wire n3258;wire n3258_t;wire WX4573;wire WX4573_t;wire n3259;wire n3259_t;wire WX4571;wire WX4571_t;wire n3260;wire n3260_t;wire WX4569;wire WX4569_t;wire n3261;wire n3261_t;wire WX4567;wire WX4567_t;wire n3262;wire n3262_t;wire WX4565;wire WX4565_t;wire n3263;wire n3263_t;wire WX4563;wire WX4563_t;wire n3264;wire n3264_t;wire WX4561;wire WX4561_t;wire n3265;wire n3265_t;wire WX4559;wire WX4559_t;wire n3266;wire n3266_t;wire WX4557;wire WX4557_t;wire n3267;wire n3267_t;wire WX4555;wire WX4555_t;wire n3268;wire n3268_t;wire WX4553;wire WX4553_t;wire WX4551;wire WX4551_t;wire WX4549;wire WX4549_t;wire WX4547;wire WX4547_t;wire WX4545;wire WX4545_t;wire WX4543;wire WX4543_t;wire WX4541;wire WX4541_t;wire WX4539;wire WX4539_t;wire WX4537;wire WX4537_t;wire WX4535;wire WX4535_t;wire WX4533;wire WX4533_t;wire WX4531;wire WX4531_t;wire WX4529;wire WX4529_t;wire WX4527;wire WX4527_t;wire WX4525;wire WX4525_t;wire WX4523;wire WX4523_t;wire WX4425;wire WX4425_t;wire WX4423;wire WX4423_t;wire WX4421;wire WX4421_t;wire WX4419;wire WX4419_t;wire WX4417;wire WX4417_t;wire WX4415;wire WX4415_t;wire WX4413;wire WX4413_t;wire WX4411;wire WX4411_t;wire WX4409;wire WX4409_t;wire WX4407;wire WX4407_t;wire WX4405;wire WX4405_t;wire WX4403;wire WX4403_t;wire WX4401;wire WX4401_t;wire WX4399;wire WX4399_t;wire WX4397;wire WX4397_t;wire WX4395;wire WX4395_t;wire WX4393;wire WX4393_t;wire WX4391;wire WX4391_t;wire WX4389;wire WX4389_t;wire WX4387;wire WX4387_t;wire WX4385;wire WX4385_t;wire WX4383;wire WX4383_t;wire WX4381;wire WX4381_t;wire WX4379;wire WX4379_t;wire WX4377;wire WX4377_t;wire WX4375;wire WX4375_t;wire WX4373;wire WX4373_t;wire WX4371;wire WX4371_t;wire WX4369;wire WX4369_t;wire WX4367;wire WX4367_t;wire WX4365;wire WX4365_t;wire WX4363;wire WX4363_t;wire WX3912;wire WX3912_t;wire WX3910;wire WX3910_t;wire WX3908;wire WX3908_t;wire WX3906;wire WX3906_t;wire WX3904;wire WX3904_t;wire WX3902;wire WX3902_t;wire WX3900;wire WX3900_t;wire WX3898;wire WX3898_t;wire WX3896;wire WX3896_t;wire WX3894;wire WX3894_t;wire WX3892;wire WX3892_t;wire WX3890;wire WX3890_t;wire WX3888;wire WX3888_t;wire WX3886;wire WX3886_t;wire WX3884;wire WX3884_t;wire WX3882;wire WX3882_t;wire WX3880;wire WX3880_t;wire WX3878;wire WX3878_t;wire WX3876;wire WX3876_t;wire WX3874;wire WX3874_t;wire WX3872;wire WX3872_t;wire WX3870;wire WX3870_t;wire WX3868;wire WX3868_t;wire WX3866;wire WX3866_t;wire WX3864;wire WX3864_t;wire WX3862;wire WX3862_t;wire WX3860;wire WX3860_t;wire WX3858;wire WX3858_t;wire WX3856;wire WX3856_t;wire WX3854;wire WX3854_t;wire WX3852;wire WX3852_t;wire WX3850;wire WX3850_t;wire WX3484;wire WX3484_t;wire WX3482;wire WX3482_t;wire WX3480;wire WX3480_t;wire WX3478;wire WX3478_t;wire WX3476;wire WX3476_t;wire WX3474;wire WX3474_t;wire WX3472;wire WX3472_t;wire WX3470;wire WX3470_t;wire WX3468;wire WX3468_t;wire WX3466;wire WX3466_t;wire WX3464;wire WX3464_t;wire WX3462;wire WX3462_t;wire WX3460;wire WX3460_t;wire WX3458;wire WX3458_t;wire WX3456;wire WX3456_t;wire WX3454;wire WX3454_t;wire WX3452;wire WX3452_t;wire WX3450;wire WX3450_t;wire WX3448;wire WX3448_t;wire WX3446;wire WX3446_t;wire WX3444;wire WX3444_t;wire WX3442;wire WX3442_t;wire WX3440;wire WX3440_t;wire WX3438;wire WX3438_t;wire WX3436;wire WX3436_t;wire WX3434;wire WX3434_t;wire WX3432;wire WX3432_t;wire WX3430;wire WX3430_t;wire WX3428;wire WX3428_t;wire WX3426;wire WX3426_t;wire WX3424;wire WX3424_t;wire WX3422;wire WX3422_t;wire WX3420;wire WX3420_t;wire WX3418;wire WX3418_t;wire WX3416;wire WX3416_t;wire WX3414;wire WX3414_t;wire WX3412;wire WX3412_t;wire WX3410;wire WX3410_t;wire WX3408;wire WX3408_t;wire WX3406;wire WX3406_t;wire WX3404;wire WX3404_t;wire WX3402;wire WX3402_t;wire WX3400;wire WX3400_t;wire WX3398;wire WX3398_t;wire WX3396;wire WX3396_t;wire WX3394;wire WX3394_t;wire WX3392;wire WX3392_t;wire WX3390;wire WX3390_t;wire WX3388;wire WX3388_t;wire WX3386;wire WX3386_t;wire WX3384;wire WX3384_t;wire WX3382;wire WX3382_t;wire WX3380;wire WX3380_t;wire WX3378;wire WX3378_t;wire WX3376;wire WX3376_t;wire WX3374;wire WX3374_t;wire WX3372;wire WX3372_t;wire WX3370;wire WX3370_t;wire WX3368;wire WX3368_t;wire WX3366;wire WX3366_t;wire WX3364;wire WX3364_t;wire WX3362;wire WX3362_t;wire WX3360;wire WX3360_t;wire WX3358;wire WX3358_t;wire WX3356;wire WX3356_t;wire WX3354;wire WX3354_t;wire WX3352;wire WX3352_t;wire WX3350;wire WX3350_t;wire WX3348;wire WX3348_t;wire WX3346;wire WX3346_t;wire WX3344;wire WX3344_t;wire WX3342;wire WX3342_t;wire WX3340;wire WX3340_t;wire WX3338;wire WX3338_t;wire WX3336;wire WX3336_t;wire WX3334;wire WX3334_t;wire WX3332;wire WX3332_t;wire WX3330;wire WX3330_t;wire WX3328;wire WX3328_t;wire WX3326;wire WX3326_t;wire WX3324;wire WX3324_t;wire WX3322;wire WX3322_t;wire WX3320;wire WX3320_t;wire WX3318;wire WX3318_t;wire WX3316;wire WX3316_t;wire WX3314;wire WX3314_t;wire WX3312;wire WX3312_t;wire WX3310;wire WX3310_t;wire WX3308;wire WX3308_t;wire WX3306;wire WX3306_t;wire WX3304;wire WX3304_t;wire WX3302;wire WX3302_t;wire WX3300;wire WX3300_t;wire WX3298;wire WX3298_t;wire WX3296;wire WX3296_t;wire WX3294;wire WX3294_t;wire WX3292;wire WX3292_t;wire n3269;wire n3269_t;wire WX3290;wire WX3290_t;wire n3270;wire n3270_t;wire WX3288;wire WX3288_t;wire n3271;wire n3271_t;wire WX3286;wire WX3286_t;wire n3272;wire n3272_t;wire WX3284;wire WX3284_t;wire n3273;wire n3273_t;wire WX3282;wire WX3282_t;wire n3274;wire n3274_t;wire WX3280;wire WX3280_t;wire n3275;wire n3275_t;wire WX3278;wire WX3278_t;wire n3276;wire n3276_t;wire WX3276;wire WX3276_t;wire n3277;wire n3277_t;wire WX3274;wire WX3274_t;wire n3278;wire n3278_t;wire WX3272;wire WX3272_t;wire n3279;wire n3279_t;wire WX3270;wire WX3270_t;wire n3280;wire n3280_t;wire WX3268;wire WX3268_t;wire n3281;wire n3281_t;wire WX3266;wire WX3266_t;wire n3282;wire n3282_t;wire WX3264;wire WX3264_t;wire n3283;wire n3283_t;wire WX3262;wire WX3262_t;wire n3284;wire n3284_t;wire WX3260;wire WX3260_t;wire WX3258;wire WX3258_t;wire WX3256;wire WX3256_t;wire WX3254;wire WX3254_t;wire WX3252;wire WX3252_t;wire WX3250;wire WX3250_t;wire WX3248;wire WX3248_t;wire WX3246;wire WX3246_t;wire WX3244;wire WX3244_t;wire WX3242;wire WX3242_t;wire WX3240;wire WX3240_t;wire WX3238;wire WX3238_t;wire WX3236;wire WX3236_t;wire WX3234;wire WX3234_t;wire WX3232;wire WX3232_t;wire WX3230;wire WX3230_t;wire WX3132;wire WX3132_t;wire WX3130;wire WX3130_t;wire WX3128;wire WX3128_t;wire WX3126;wire WX3126_t;wire WX3124;wire WX3124_t;wire WX3122;wire WX3122_t;wire WX3120;wire WX3120_t;wire WX3118;wire WX3118_t;wire WX3116;wire WX3116_t;wire WX3114;wire WX3114_t;wire WX3112;wire WX3112_t;wire WX3110;wire WX3110_t;wire WX3108;wire WX3108_t;wire WX3106;wire WX3106_t;wire WX3104;wire WX3104_t;wire WX3102;wire WX3102_t;wire WX3100;wire WX3100_t;wire WX3098;wire WX3098_t;wire WX3096;wire WX3096_t;wire WX3094;wire WX3094_t;wire WX3092;wire WX3092_t;wire WX3090;wire WX3090_t;wire WX3088;wire WX3088_t;wire WX3086;wire WX3086_t;wire WX3084;wire WX3084_t;wire WX3082;wire WX3082_t;wire WX3080;wire WX3080_t;wire WX3078;wire WX3078_t;wire WX3076;wire WX3076_t;wire WX3074;wire WX3074_t;wire WX3072;wire WX3072_t;wire WX3070;wire WX3070_t;wire WX2619;wire WX2619_t;wire WX2617;wire WX2617_t;wire WX2615;wire WX2615_t;wire WX2613;wire WX2613_t;wire WX2611;wire WX2611_t;wire WX2609;wire WX2609_t;wire WX2607;wire WX2607_t;wire WX2605;wire WX2605_t;wire WX2603;wire WX2603_t;wire WX2601;wire WX2601_t;wire WX2599;wire WX2599_t;wire WX2597;wire WX2597_t;wire WX2595;wire WX2595_t;wire WX2593;wire WX2593_t;wire WX2591;wire WX2591_t;wire WX2589;wire WX2589_t;wire WX2587;wire WX2587_t;wire WX2585;wire WX2585_t;wire WX2583;wire WX2583_t;wire WX2581;wire WX2581_t;wire WX2579;wire WX2579_t;wire WX2577;wire WX2577_t;wire WX2575;wire WX2575_t;wire WX2573;wire WX2573_t;wire WX2571;wire WX2571_t;wire WX2569;wire WX2569_t;wire WX2567;wire WX2567_t;wire WX2565;wire WX2565_t;wire WX2563;wire WX2563_t;wire WX2561;wire WX2561_t;wire WX2559;wire WX2559_t;wire WX2557;wire WX2557_t;wire WX2191;wire WX2191_t;wire WX2189;wire WX2189_t;wire WX2187;wire WX2187_t;wire WX2185;wire WX2185_t;wire WX2183;wire WX2183_t;wire WX2181;wire WX2181_t;wire WX2179;wire WX2179_t;wire WX2177;wire WX2177_t;wire WX2175;wire WX2175_t;wire WX2173;wire WX2173_t;wire WX2171;wire WX2171_t;wire WX2169;wire WX2169_t;wire WX2167;wire WX2167_t;wire WX2165;wire WX2165_t;wire WX2163;wire WX2163_t;wire WX2161;wire WX2161_t;wire WX2159;wire WX2159_t;wire WX2157;wire WX2157_t;wire WX2155;wire WX2155_t;wire WX2153;wire WX2153_t;wire WX2151;wire WX2151_t;wire WX2149;wire WX2149_t;wire WX2147;wire WX2147_t;wire WX2145;wire WX2145_t;wire WX2143;wire WX2143_t;wire WX2141;wire WX2141_t;wire WX2139;wire WX2139_t;wire WX2137;wire WX2137_t;wire WX2135;wire WX2135_t;wire WX2133;wire WX2133_t;wire WX2131;wire WX2131_t;wire WX2129;wire WX2129_t;wire WX2127;wire WX2127_t;wire WX2125;wire WX2125_t;wire WX2123;wire WX2123_t;wire WX2121;wire WX2121_t;wire WX2119;wire WX2119_t;wire WX2117;wire WX2117_t;wire WX2115;wire WX2115_t;wire WX2113;wire WX2113_t;wire WX2111;wire WX2111_t;wire WX2109;wire WX2109_t;wire WX2107;wire WX2107_t;wire WX2105;wire WX2105_t;wire WX2103;wire WX2103_t;wire WX2101;wire WX2101_t;wire WX2099;wire WX2099_t;wire WX2097;wire WX2097_t;wire WX2095;wire WX2095_t;wire WX2093;wire WX2093_t;wire WX2091;wire WX2091_t;wire WX2089;wire WX2089_t;wire WX2087;wire WX2087_t;wire WX2085;wire WX2085_t;wire WX2083;wire WX2083_t;wire WX2081;wire WX2081_t;wire WX2079;wire WX2079_t;wire WX2077;wire WX2077_t;wire WX2075;wire WX2075_t;wire WX2073;wire WX2073_t;wire WX2071;wire WX2071_t;wire WX2069;wire WX2069_t;wire WX2067;wire WX2067_t;wire WX2065;wire WX2065_t;wire WX2063;wire WX2063_t;wire WX2061;wire WX2061_t;wire WX2059;wire WX2059_t;wire WX2057;wire WX2057_t;wire WX2055;wire WX2055_t;wire WX2053;wire WX2053_t;wire WX2051;wire WX2051_t;wire WX2049;wire WX2049_t;wire WX2047;wire WX2047_t;wire WX2045;wire WX2045_t;wire WX2043;wire WX2043_t;wire WX2041;wire WX2041_t;wire WX2039;wire WX2039_t;wire WX2037;wire WX2037_t;wire WX2035;wire WX2035_t;wire WX2033;wire WX2033_t;wire WX2031;wire WX2031_t;wire WX2029;wire WX2029_t;wire WX2027;wire WX2027_t;wire WX2025;wire WX2025_t;wire WX2023;wire WX2023_t;wire WX2021;wire WX2021_t;wire WX2019;wire WX2019_t;wire WX2017;wire WX2017_t;wire WX2015;wire WX2015_t;wire WX2013;wire WX2013_t;wire WX2011;wire WX2011_t;wire WX2009;wire WX2009_t;wire WX2007;wire WX2007_t;wire WX2005;wire WX2005_t;wire WX2003;wire WX2003_t;wire WX2001;wire WX2001_t;wire WX1999;wire WX1999_t;wire n3285;wire n3285_t;wire n3286;wire n3286_t;wire WX1997;wire WX1997_t;wire n3287;wire n3287_t;wire n3288;wire n3288_t;wire WX1995;wire WX1995_t;wire n3289;wire n3289_t;wire n3290;wire n3290_t;wire WX1993;wire WX1993_t;wire n3291;wire n3291_t;wire n3292;wire n3292_t;wire WX1991;wire WX1991_t;wire n3293;wire n3293_t;wire n3294;wire n3294_t;wire WX1989;wire WX1989_t;wire n3295;wire n3295_t;wire n3296;wire n3296_t;wire WX1987;wire WX1987_t;wire n3297;wire n3297_t;wire n3298;wire n3298_t;wire WX1985;wire WX1985_t;wire n3299;wire n3299_t;wire n3300;wire n3300_t;wire WX1983;wire WX1983_t;wire n3301;wire n3301_t;wire n3302;wire n3302_t;wire WX1981;wire WX1981_t;wire n3303;wire n3303_t;wire n3304;wire n3304_t;wire WX1979;wire WX1979_t;wire n3305;wire n3305_t;wire n3306;wire n3306_t;wire WX1977;wire WX1977_t;wire n3307;wire n3307_t;wire n3308;wire n3308_t;wire WX1975;wire WX1975_t;wire n3309;wire n3309_t;wire n3310;wire n3310_t;wire WX1973;wire WX1973_t;wire n3311;wire n3311_t;wire n3312;wire n3312_t;wire WX1971;wire WX1971_t;wire n3313;wire n3313_t;wire n3314;wire n3314_t;wire WX1969;wire WX1969_t;wire n3315;wire n3315_t;wire n3316;wire n3316_t;wire WX1967;wire WX1967_t;wire WX1965;wire WX1965_t;wire WX1963;wire WX1963_t;wire WX1961;wire WX1961_t;wire WX1959;wire WX1959_t;wire WX1957;wire WX1957_t;wire WX1955;wire WX1955_t;wire WX1953;wire WX1953_t;wire WX1951;wire WX1951_t;wire WX1949;wire WX1949_t;wire WX1947;wire WX1947_t;wire WX1945;wire WX1945_t;wire WX1943;wire WX1943_t;wire WX1941;wire WX1941_t;wire WX1939;wire WX1939_t;wire WX1937;wire WX1937_t;wire WX1839;wire WX1839_t;wire WX1837;wire WX1837_t;wire WX1835;wire WX1835_t;wire WX1833;wire WX1833_t;wire WX1831;wire WX1831_t;wire WX1829;wire WX1829_t;wire WX1827;wire WX1827_t;wire WX1825;wire WX1825_t;wire WX1823;wire WX1823_t;wire WX1821;wire WX1821_t;wire WX1819;wire WX1819_t;wire WX1817;wire WX1817_t;wire WX1815;wire WX1815_t;wire WX1813;wire WX1813_t;wire WX1811;wire WX1811_t;wire WX1809;wire WX1809_t;wire WX1807;wire WX1807_t;wire WX1805;wire WX1805_t;wire WX1803;wire WX1803_t;wire WX1801;wire WX1801_t;wire WX1799;wire WX1799_t;wire WX1797;wire WX1797_t;wire WX1795;wire WX1795_t;wire WX1793;wire WX1793_t;wire WX1791;wire WX1791_t;wire WX1789;wire WX1789_t;wire WX1787;wire WX1787_t;wire WX1785;wire WX1785_t;wire WX1783;wire WX1783_t;wire WX1781;wire WX1781_t;wire WX1779;wire WX1779_t;wire WX1777;wire WX1777_t;wire WX1326;wire WX1326_t;wire WX1324;wire WX1324_t;wire WX1322;wire WX1322_t;wire WX1320;wire WX1320_t;wire WX1318;wire WX1318_t;wire WX1316;wire WX1316_t;wire WX1314;wire WX1314_t;wire WX1312;wire WX1312_t;wire WX1310;wire WX1310_t;wire WX1308;wire WX1308_t;wire WX1306;wire WX1306_t;wire WX1304;wire WX1304_t;wire WX1302;wire WX1302_t;wire WX1300;wire WX1300_t;wire WX1298;wire WX1298_t;wire WX1296;wire WX1296_t;wire WX1294;wire WX1294_t;wire WX1292;wire WX1292_t;wire WX1290;wire WX1290_t;wire WX1288;wire WX1288_t;wire WX1286;wire WX1286_t;wire WX1284;wire WX1284_t;wire WX1282;wire WX1282_t;wire WX1280;wire WX1280_t;wire WX1278;wire WX1278_t;wire WX1276;wire WX1276_t;wire WX1274;wire WX1274_t;wire WX1272;wire WX1272_t;wire WX1270;wire WX1270_t;wire WX1268;wire WX1268_t;wire WX1266;wire WX1266_t;wire WX1264;wire WX1264_t;wire WX11670;wire WX11670_t;wire WX11668;wire WX11668_t;wire WX11666;wire WX11666_t;wire WX11664;wire WX11664_t;wire WX11662;wire WX11662_t;wire WX11660;wire WX11660_t;wire WX11658;wire WX11658_t;wire WX11656;wire WX11656_t;wire WX11654;wire WX11654_t;wire WX11652;wire WX11652_t;wire WX11650;wire WX11650_t;wire WX11648;wire WX11648_t;wire WX11646;wire WX11646_t;wire WX11644;wire WX11644_t;wire WX11642;wire WX11642_t;wire WX11640;wire WX11640_t;wire WX11638;wire WX11638_t;wire WX11636;wire WX11636_t;wire WX11634;wire WX11634_t;wire WX11632;wire WX11632_t;wire WX11630;wire WX11630_t;wire WX11628;wire WX11628_t;wire WX11626;wire WX11626_t;wire WX11624;wire WX11624_t;wire WX11622;wire WX11622_t;wire WX11620;wire WX11620_t;wire WX11618;wire WX11618_t;wire WX11616;wire WX11616_t;wire WX11614;wire WX11614_t;wire WX11612;wire WX11612_t;wire WX11610;wire WX11610_t;wire WX11608;wire WX11608_t;wire WX11242;wire WX11242_t;wire WX11240;wire WX11240_t;wire WX11238;wire WX11238_t;wire WX11236;wire WX11236_t;wire WX11234;wire WX11234_t;wire WX11232;wire WX11232_t;wire WX11230;wire WX11230_t;wire WX11228;wire WX11228_t;wire WX11226;wire WX11226_t;wire WX11224;wire WX11224_t;wire WX11222;wire WX11222_t;wire WX11220;wire WX11220_t;wire WX11218;wire WX11218_t;wire WX11216;wire WX11216_t;wire WX11214;wire WX11214_t;wire WX11212;wire WX11212_t;wire WX11210;wire WX11210_t;wire WX11208;wire WX11208_t;wire WX11206;wire WX11206_t;wire WX11204;wire WX11204_t;wire WX11202;wire WX11202_t;wire WX11200;wire WX11200_t;wire WX11198;wire WX11198_t;wire WX11196;wire WX11196_t;wire WX11194;wire WX11194_t;wire WX11192;wire WX11192_t;wire WX11190;wire WX11190_t;wire WX11188;wire WX11188_t;wire WX11186;wire WX11186_t;wire WX11184;wire WX11184_t;wire WX11182;wire WX11182_t;wire WX11180;wire WX11180_t;wire WX11178;wire WX11178_t;wire WX11176;wire WX11176_t;wire WX11174;wire WX11174_t;wire WX11172;wire WX11172_t;wire WX11170;wire WX11170_t;wire WX11168;wire WX11168_t;wire WX11166;wire WX11166_t;wire WX11164;wire WX11164_t;wire WX11162;wire WX11162_t;wire WX11160;wire WX11160_t;wire WX11158;wire WX11158_t;wire WX11156;wire WX11156_t;wire WX11154;wire WX11154_t;wire WX11152;wire WX11152_t;wire WX11150;wire WX11150_t;wire WX11148;wire WX11148_t;wire WX11146;wire WX11146_t;wire WX11144;wire WX11144_t;wire WX11142;wire WX11142_t;wire WX11140;wire WX11140_t;wire WX11138;wire WX11138_t;wire WX11136;wire WX11136_t;wire WX11134;wire WX11134_t;wire WX11132;wire WX11132_t;wire WX11130;wire WX11130_t;wire WX11128;wire WX11128_t;wire WX11126;wire WX11126_t;wire WX11124;wire WX11124_t;wire WX11122;wire WX11122_t;wire WX11120;wire WX11120_t;wire WX11118;wire WX11118_t;wire WX11116;wire WX11116_t;wire WX11114;wire WX11114_t;wire WX11112;wire WX11112_t;wire WX11110;wire WX11110_t;wire WX11108;wire WX11108_t;wire WX11106;wire WX11106_t;wire WX11104;wire WX11104_t;wire WX11102;wire WX11102_t;wire WX11100;wire WX11100_t;wire WX11098;wire WX11098_t;wire WX11096;wire WX11096_t;wire WX11094;wire WX11094_t;wire WX11092;wire WX11092_t;wire WX11090;wire WX11090_t;wire WX11088;wire WX11088_t;wire WX11086;wire WX11086_t;wire WX11084;wire WX11084_t;wire WX11082;wire WX11082_t;wire WX11080;wire WX11080_t;wire WX11078;wire WX11078_t;wire WX11076;wire WX11076_t;wire WX11074;wire WX11074_t;wire WX11072;wire WX11072_t;wire WX11070;wire WX11070_t;wire WX11068;wire WX11068_t;wire WX11066;wire WX11066_t;wire WX11064;wire WX11064_t;wire WX11062;wire WX11062_t;wire WX11060;wire WX11060_t;wire WX11058;wire WX11058_t;wire WX11056;wire WX11056_t;wire WX11054;wire WX11054_t;wire WX11052;wire WX11052_t;wire WX11050;wire WX11050_t;wire n3317;wire n3317_t;wire WX11048;wire WX11048_t;wire n3318;wire n3318_t;wire WX11046;wire WX11046_t;wire n3319;wire n3319_t;wire WX11044;wire WX11044_t;wire n3320;wire n3320_t;wire WX11042;wire WX11042_t;wire n3321;wire n3321_t;wire WX11040;wire WX11040_t;wire n3322;wire n3322_t;wire WX11038;wire WX11038_t;wire n3323;wire n3323_t;wire WX11036;wire WX11036_t;wire n3324;wire n3324_t;wire WX11034;wire WX11034_t;wire n3325;wire n3325_t;wire WX11032;wire WX11032_t;wire n3326;wire n3326_t;wire WX11030;wire WX11030_t;wire n3327;wire n3327_t;wire WX11028;wire WX11028_t;wire n3328;wire n3328_t;wire WX11026;wire WX11026_t;wire n3329;wire n3329_t;wire WX11024;wire WX11024_t;wire n3330;wire n3330_t;wire WX11022;wire WX11022_t;wire n3331;wire n3331_t;wire WX11020;wire WX11020_t;wire n3332;wire n3332_t;wire WX11018;wire WX11018_t;wire WX11016;wire WX11016_t;wire WX11014;wire WX11014_t;wire WX11012;wire WX11012_t;wire WX11010;wire WX11010_t;wire WX11008;wire WX11008_t;wire WX11006;wire WX11006_t;wire WX11004;wire WX11004_t;wire WX11002;wire WX11002_t;wire WX11000;wire WX11000_t;wire WX10998;wire WX10998_t;wire WX10996;wire WX10996_t;wire WX10994;wire WX10994_t;wire WX10992;wire WX10992_t;wire WX10990;wire WX10990_t;wire WX10988;wire WX10988_t;wire WX10890;wire WX10890_t;wire WX10888;wire WX10888_t;wire WX10886;wire WX10886_t;wire WX10884;wire WX10884_t;wire WX10882;wire WX10882_t;wire WX10880;wire WX10880_t;wire WX10878;wire WX10878_t;wire WX10876;wire WX10876_t;wire WX10874;wire WX10874_t;wire WX10872;wire WX10872_t;wire WX10870;wire WX10870_t;wire WX10868;wire WX10868_t;wire WX10866;wire WX10866_t;wire WX10864;wire WX10864_t;wire WX10862;wire WX10862_t;wire WX10860;wire WX10860_t;wire WX10858;wire WX10858_t;wire WX10856;wire WX10856_t;wire WX10854;wire WX10854_t;wire WX10852;wire WX10852_t;wire WX10850;wire WX10850_t;wire WX10848;wire WX10848_t;wire WX10846;wire WX10846_t;wire WX10844;wire WX10844_t;wire WX10842;wire WX10842_t;wire WX10840;wire WX10840_t;wire WX10838;wire WX10838_t;wire WX10836;wire WX10836_t;wire WX10834;wire WX10834_t;wire WX10832;wire WX10832_t;wire WX10830;wire WX10830_t;wire WX10828;wire WX10828_t;wire WX10377;wire WX10377_t;wire WX10375;wire WX10375_t;wire WX10373;wire WX10373_t;wire WX10371;wire WX10371_t;wire WX10369;wire WX10369_t;wire WX10367;wire WX10367_t;wire WX10365;wire WX10365_t;wire WX10363;wire WX10363_t;wire WX10361;wire WX10361_t;wire WX10359;wire WX10359_t;wire WX10357;wire WX10357_t;wire WX10355;wire WX10355_t;wire WX10353;wire WX10353_t;wire WX10351;wire WX10351_t;wire WX10349;wire WX10349_t;wire WX10347;wire WX10347_t;wire WX10345;wire WX10345_t;wire WX10343;wire WX10343_t;wire WX10341;wire WX10341_t;wire WX10339;wire WX10339_t;wire WX10337;wire WX10337_t;wire WX10335;wire WX10335_t;wire WX10333;wire WX10333_t;wire WX10331;wire WX10331_t;wire WX10329;wire WX10329_t;wire WX10327;wire WX10327_t;wire WX10325;wire WX10325_t;wire WX10323;wire WX10323_t;wire WX10321;wire WX10321_t;wire WX10319;wire WX10319_t;wire WX10317;wire WX10317_t;wire WX10315;wire WX10315_t;wire n1729;wire n1729_t;wire n1730;wire n1730_t;wire n1731;wire n1731_t;wire n1732;wire n1732_t;wire n1733;wire n1733_t;wire n1734;wire n1734_t;wire n1735;wire n1735_t;wire n1736;wire n1736_t;wire n1737;wire n1737_t;wire n1738;wire n1738_t;wire n1739;wire n1739_t;wire n1740;wire n1740_t;wire n1741;wire n1741_t;wire n1742;wire n1742_t;wire n1743;wire n1743_t;wire n1744;wire n1744_t;wire n1745;wire n1745_t;wire n1746;wire n1746_t;wire n1747;wire n1747_t;wire n1748;wire n1748_t;wire n1749;wire n1749_t;wire n1750;wire n1750_t;wire n1751;wire n1751_t;wire n1752;wire n1752_t;wire n1753;wire n1753_t;wire n1754;wire n1754_t;wire n1755;wire n1755_t;wire n1756;wire n1756_t;wire n1757;wire n1757_t;wire n1758;wire n1758_t;wire n1759;wire n1759_t;wire n1760;wire n1760_t;wire n1761;wire n1761_t;wire n1762;wire n1762_t;wire n1763;wire n1763_t;wire n1764;wire n1764_t;wire n1765;wire n1765_t;wire n1766;wire n1766_t;wire n1767;wire n1767_t;wire n1768;wire n1768_t;wire n1769;wire n1769_t;wire n1770;wire n1770_t;wire n1771;wire n1771_t;wire n1772;wire n1772_t;wire n1773;wire n1773_t;wire n1774;wire n1774_t;wire n1775;wire n1775_t;wire n1776;wire n1776_t;wire n1777;wire n1777_t;wire n1778;wire n1778_t;wire n1779;wire n1779_t;wire n1780;wire n1780_t;wire n1781;wire n1781_t;wire n1782;wire n1782_t;wire n1783;wire n1783_t;wire n1784;wire n1784_t;wire n1785;wire n1785_t;wire n1786;wire n1786_t;wire n1787;wire n1787_t;wire n1788;wire n1788_t;wire n1789;wire n1789_t;wire n1790;wire n1790_t;wire n1791;wire n1791_t;wire n1792;wire n1792_t;wire n1793;wire n1793_t;wire n1794;wire n1794_t;wire n1795;wire n1795_t;wire n1796;wire n1796_t;wire n1797;wire n1797_t;wire n1798;wire n1798_t;wire n1799;wire n1799_t;wire n1800;wire n1800_t;wire n1801;wire n1801_t;wire n1802;wire n1802_t;wire n1803;wire n1803_t;wire n1804;wire n1804_t;wire n1805;wire n1805_t;wire n1806;wire n1806_t;wire n1807;wire n1807_t;wire n1808;wire n1808_t;wire n1809;wire n1809_t;wire n1810;wire n1810_t;wire n1811;wire n1811_t;wire n1812;wire n1812_t;wire n1813;wire n1813_t;wire n1814;wire n1814_t;wire n1815;wire n1815_t;wire n1816;wire n1816_t;wire n1817;wire n1817_t;wire n1818;wire n1818_t;wire n1819;wire n1819_t;wire n1820;wire n1820_t;wire n1821;wire n1821_t;wire n1822;wire n1822_t;wire n1823;wire n1823_t;wire n1824;wire n1824_t;wire n1825;wire n1825_t;wire n1826;wire n1826_t;wire n1827;wire n1827_t;wire n1828;wire n1828_t;wire n1829;wire n1829_t;wire n1830;wire n1830_t;wire n1831;wire n1831_t;wire n1832;wire n1832_t;wire n1833;wire n1833_t;wire n1834;wire n1834_t;wire n1835;wire n1835_t;wire n1836;wire n1836_t;wire n1837;wire n1837_t;wire n1838;wire n1838_t;wire n1839;wire n1839_t;wire n1840;wire n1840_t;wire n1841;wire n1841_t;wire n1842;wire n1842_t;wire n1843;wire n1843_t;wire n1844;wire n1844_t;wire n1845;wire n1845_t;wire n1846;wire n1846_t;wire n1847;wire n1847_t;wire n1848;wire n1848_t;wire n1849;wire n1849_t;wire n1850;wire n1850_t;wire n1851;wire n1851_t;wire n1852;wire n1852_t;wire n1853;wire n1853_t;wire n1854;wire n1854_t;wire n1855;wire n1855_t;wire n1856;wire n1856_t;wire n1857;wire n1857_t;wire n1858;wire n1858_t;wire n1859;wire n1859_t;wire n1860;wire n1860_t;wire n1861;wire n1861_t;wire n1862;wire n1862_t;wire n1863;wire n1863_t;wire n1864;wire n1864_t;wire n1865;wire n1865_t;wire n1866;wire n1866_t;wire n1867;wire n1867_t;wire n1868;wire n1868_t;wire n1869;wire n1869_t;wire n1870;wire n1870_t;wire n1871;wire n1871_t;wire n1872;wire n1872_t;wire n1873;wire n1873_t;wire n1874;wire n1874_t;wire n1875;wire n1875_t;wire n1876;wire n1876_t;wire n1877;wire n1877_t;wire n1878;wire n1878_t;wire n1879;wire n1879_t;wire n1880;wire n1880_t;wire n1881;wire n1881_t;wire n1882;wire n1882_t;wire n1883;wire n1883_t;wire n1884;wire n1884_t;wire n1885;wire n1885_t;wire n1886;wire n1886_t;wire n1887;wire n1887_t;wire n1888;wire n1888_t;wire n1889;wire n1889_t;wire n1890;wire n1890_t;wire n1891;wire n1891_t;wire n1892;wire n1892_t;wire n1893;wire n1893_t;wire n1894;wire n1894_t;wire n1895;wire n1895_t;wire n1896;wire n1896_t;wire n1897;wire n1897_t;wire n1898;wire n1898_t;wire n1899;wire n1899_t;wire n1900;wire n1900_t;wire n1901;wire n1901_t;wire n1902;wire n1902_t;wire n1903;wire n1903_t;wire n1904;wire n1904_t;wire n1905;wire n1905_t;wire n1906;wire n1906_t;wire n1907;wire n1907_t;wire n1908;wire n1908_t;wire n1909;wire n1909_t;wire n1910;wire n1910_t;wire n1911;wire n1911_t;wire n1912;wire n1912_t;wire n1913;wire n1913_t;wire n1914;wire n1914_t;wire n1915;wire n1915_t;wire n1916;wire n1916_t;wire n1917;wire n1917_t;wire n1918;wire n1918_t;wire n1919;wire n1919_t;wire n1920;wire n1920_t;wire n1921;wire n1921_t;wire n1922;wire n1922_t;wire n1923;wire n1923_t;wire n1924;wire n1924_t;wire n1925;wire n1925_t;wire n1926;wire n1926_t;wire n1927;wire n1927_t;wire n1928;wire n1928_t;wire n1929;wire n1929_t;wire n1930;wire n1930_t;wire n1931;wire n1931_t;wire n1932;wire n1932_t;wire n1933;wire n1933_t;wire n1934;wire n1934_t;wire n1935;wire n1935_t;wire n1936;wire n1936_t;wire n1937;wire n1937_t;wire n1938;wire n1938_t;wire n1939;wire n1939_t;wire n1940;wire n1940_t;wire n1941;wire n1941_t;wire n1942;wire n1942_t;wire n1943;wire n1943_t;wire n1944;wire n1944_t;wire n1945;wire n1945_t;wire n1946;wire n1946_t;wire n1947;wire n1947_t;wire n1948;wire n1948_t;wire n1949;wire n1949_t;wire n1950;wire n1950_t;wire n1951;wire n1951_t;wire n1952;wire n1952_t;wire n1953;wire n1953_t;wire n1954;wire n1954_t;wire n1955;wire n1955_t;wire n1956;wire n1956_t;wire n1957;wire n1957_t;wire n1958;wire n1958_t;wire n1959;wire n1959_t;wire n1960;wire n1960_t;wire n1961;wire n1961_t;wire n1962;wire n1962_t;wire n1963;wire n1963_t;wire n1964;wire n1964_t;wire n1965;wire n1965_t;wire n1966;wire n1966_t;wire n1967;wire n1967_t;wire n1968;wire n1968_t;wire n1969;wire n1969_t;wire n1970;wire n1970_t;wire n1971;wire n1971_t;wire n1972;wire n1972_t;wire n1973;wire n1973_t;wire n1974;wire n1974_t;wire n1975;wire n1975_t;wire n1976;wire n1976_t;wire n1977;wire n1977_t;wire n1978;wire n1978_t;wire n1979;wire n1979_t;wire n1980;wire n1980_t;wire n1981;wire n1981_t;wire n1982;wire n1982_t;wire n1983;wire n1983_t;wire n1984;wire n1984_t;wire n1985;wire n1985_t;wire n1986;wire n1986_t;wire n1987;wire n1987_t;wire n1988;wire n1988_t;wire n1989;wire n1989_t;wire n1990;wire n1990_t;wire n1991;wire n1991_t;wire n1992;wire n1992_t;wire n1993;wire n1993_t;wire n1994;wire n1994_t;wire n1995;wire n1995_t;wire n1996;wire n1996_t;wire n1997;wire n1997_t;wire n1998;wire n1998_t;wire n1999;wire n1999_t;wire n2000;wire n2000_t;wire n2001;wire n2001_t;wire n2002;wire n2002_t;wire n2003;wire n2003_t;wire n2004;wire n2004_t;wire n2005;wire n2005_t;wire n2006;wire n2006_t;wire n2007;wire n2007_t;wire n2008;wire n2008_t;wire n2009;wire n2009_t;wire n2010;wire n2010_t;wire n2011;wire n2011_t;wire n2012;wire n2012_t;wire n2013;wire n2013_t;wire n2014;wire n2014_t;wire n2015;wire n2015_t;wire n2016;wire n2016_t;wire n2017;wire n2017_t;wire n2018;wire n2018_t;wire n2019;wire n2019_t;wire n2020;wire n2020_t;wire n2021;wire n2021_t;wire n2022;wire n2022_t;wire n2023;wire n2023_t;wire n2024;wire n2024_t;wire n2025;wire n2025_t;wire n2026;wire n2026_t;wire n2027;wire n2027_t;wire n2028;wire n2028_t;wire n2029;wire n2029_t;wire n2030;wire n2030_t;wire n2031;wire n2031_t;wire n2032;wire n2032_t;wire n2033;wire n2033_t;wire n2034;wire n2034_t;wire n2035;wire n2035_t;wire n2036;wire n2036_t;wire n2037;wire n2037_t;wire n2038;wire n2038_t;wire n2039;wire n2039_t;wire n2040;wire n2040_t;wire n2041;wire n2041_t;wire n2042;wire n2042_t;wire n2043;wire n2043_t;wire n2044;wire n2044_t;wire n2045;wire n2045_t;wire n2046;wire n2046_t;wire n2047;wire n2047_t;wire n2048;wire n2048_t;wire n2049;wire n2049_t;wire n2050;wire n2050_t;wire n2051;wire n2051_t;wire n2052;wire n2052_t;wire n2053;wire n2053_t;wire n2054;wire n2054_t;wire n2055;wire n2055_t;wire n2056;wire n2056_t;wire n2057;wire n2057_t;wire n2058;wire n2058_t;wire n2059;wire n2059_t;wire n2060;wire n2060_t;wire n2061;wire n2061_t;wire n2062;wire n2062_t;wire n2063;wire n2063_t;wire n2064;wire n2064_t;wire n2065;wire n2065_t;wire n2066;wire n2066_t;wire n2067;wire n2067_t;wire n2068;wire n2068_t;wire n2069;wire n2069_t;wire n2070;wire n2070_t;wire n2071;wire n2071_t;wire n2072;wire n2072_t;wire n2073;wire n2073_t;wire n2074;wire n2074_t;wire n2075;wire n2075_t;wire n2076;wire n2076_t;wire n2077;wire n2077_t;wire n2078;wire n2078_t;wire n2079;wire n2079_t;wire n2080;wire n2080_t;wire n2081;wire n2081_t;wire n2082;wire n2082_t;wire n2083;wire n2083_t;wire n2084;wire n2084_t;wire n2085;wire n2085_t;wire n2086;wire n2086_t;wire n2087;wire n2087_t;wire n2088;wire n2088_t;wire n2089;wire n2089_t;wire n2090;wire n2090_t;wire n2091;wire n2091_t;wire n2092;wire n2092_t;wire n2093;wire n2093_t;wire n2094;wire n2094_t;wire n2095;wire n2095_t;wire n2096;wire n2096_t;wire n2097;wire n2097_t;wire n2098;wire n2098_t;wire n2099;wire n2099_t;wire n2100;wire n2100_t;wire n2101;wire n2101_t;wire n2102;wire n2102_t;wire n2103;wire n2103_t;wire n2104;wire n2104_t;wire n2105;wire n2105_t;wire n2106;wire n2106_t;wire n2107;wire n2107_t;wire n2108;wire n2108_t;wire n2109;wire n2109_t;wire n2110;wire n2110_t;wire n2111;wire n2111_t;wire n2112;wire n2112_t;wire n2113;wire n2113_t;wire n2114;wire n2114_t;wire n2115;wire n2115_t;wire n2116;wire n2116_t;wire n2117;wire n2117_t;wire n2118;wire n2118_t;wire n2119;wire n2119_t;wire n2120;wire n2120_t;wire n2121;wire n2121_t;wire n2122;wire n2122_t;wire n2123;wire n2123_t;wire n2124;wire n2124_t;wire n2125;wire n2125_t;wire n2126;wire n2126_t;wire n2127;wire n2127_t;wire n2128;wire n2128_t;wire n2129;wire n2129_t;wire n2130;wire n2130_t;wire n2131;wire n2131_t;wire n2132;wire n2132_t;wire n2133;wire n2133_t;wire n2134;wire n2134_t;wire n2135;wire n2135_t;wire n2136;wire n2136_t;wire n2137;wire n2137_t;wire n2138;wire n2138_t;wire n2139;wire n2139_t;wire n2140;wire n2140_t;wire n2141;wire n2141_t;wire n2142;wire n2142_t;wire n2143;wire n2143_t;wire n2144;wire n2144_t;wire n2145;wire n2145_t;wire n2146;wire n2146_t;wire n2147;wire n2147_t;wire n2148;wire n2148_t;wire n2149;wire n2149_t;wire n2150;wire n2150_t;wire n2151;wire n2151_t;wire n2152;wire n2152_t;wire n2153;wire n2153_t;wire n2154;wire n2154_t;wire n2155;wire n2155_t;wire n2156;wire n2156_t;wire n2157;wire n2157_t;wire n2158;wire n2158_t;wire n2159;wire n2159_t;wire n2160;wire n2160_t;wire n2161;wire n2161_t;wire n2162;wire n2162_t;wire n2163;wire n2163_t;wire n2164;wire n2164_t;wire n2165;wire n2165_t;wire n2166;wire n2166_t;wire n2167;wire n2167_t;wire n2168;wire n2168_t;wire n2169;wire n2169_t;wire n2170;wire n2170_t;wire n2171;wire n2171_t;wire n2172;wire n2172_t;wire n2173;wire n2173_t;wire n2174;wire n2174_t;wire n2175;wire n2175_t;wire n2176;wire n2176_t;wire n2177;wire n2177_t;wire n2178;wire n2178_t;wire n2179;wire n2179_t;wire n2180;wire n2180_t;wire n2181;wire n2181_t;wire n2182;wire n2182_t;wire n2183;wire n2183_t;wire n2184;wire n2184_t;wire n2185;wire n2185_t;wire n2186;wire n2186_t;wire n2187;wire n2187_t;wire n2188;wire n2188_t;wire n2189;wire n2189_t;wire n2190;wire n2190_t;wire n2191;wire n2191_t;wire n2192;wire n2192_t;wire n2193;wire n2193_t;wire n2194;wire n2194_t;wire n2195;wire n2195_t;wire n2196;wire n2196_t;wire n2197;wire n2197_t;wire n2198;wire n2198_t;wire n2199;wire n2199_t;wire n2200;wire n2200_t;wire n2201;wire n2201_t;wire n2202;wire n2202_t;wire n2203;wire n2203_t;wire n2204;wire n2204_t;wire n2205;wire n2205_t;wire n2206;wire n2206_t;wire n2207;wire n2207_t;wire n2208;wire n2208_t;wire n2209;wire n2209_t;wire n2210;wire n2210_t;wire n2211;wire n2211_t;wire n2212;wire n2212_t;wire n2213;wire n2213_t;wire n2214;wire n2214_t;wire n2215;wire n2215_t;wire n2216;wire n2216_t;wire n2217;wire n2217_t;wire n2218;wire n2218_t;wire n2219;wire n2219_t;wire n2220;wire n2220_t;wire n2221;wire n2221_t;wire n2222;wire n2222_t;wire n2223;wire n2223_t;wire n2224;wire n2224_t;wire n2225;wire n2225_t;wire n2226;wire n2226_t;wire n2227;wire n2227_t;wire n2228;wire n2228_t;wire n2229;wire n2229_t;wire n2230;wire n2230_t;wire n2231;wire n2231_t;wire n2232;wire n2232_t;wire n2233;wire n2233_t;wire n2234;wire n2234_t;wire n2235;wire n2235_t;wire n2236;wire n2236_t;wire n2237;wire n2237_t;wire n2238;wire n2238_t;wire n2239;wire n2239_t;wire n2240;wire n2240_t;wire n2241;wire n2241_t;wire n2242;wire n2242_t;wire n2243;wire n2243_t;wire n2244;wire n2244_t;wire n2245;wire n2245_t;wire n2246;wire n2246_t;wire n2247;wire n2247_t;wire n2248;wire n2248_t;wire n2249;wire n2249_t;wire n2250;wire n2250_t;wire n2251;wire n2251_t;wire n2252;wire n2252_t;wire n2253;wire n2253_t;wire n2254;wire n2254_t;wire n2255;wire n2255_t;wire n2256;wire n2256_t;wire n2257;wire n2257_t;wire n2258;wire n2258_t;wire n2259;wire n2259_t;wire n2260;wire n2260_t;wire n2261;wire n2261_t;wire n2262;wire n2262_t;wire n2263;wire n2263_t;wire n2264;wire n2264_t;wire n2265;wire n2265_t;wire n2266;wire n2266_t;wire n2267;wire n2267_t;wire n2268;wire n2268_t;wire n2269;wire n2269_t;wire n2270;wire n2270_t;wire n2271;wire n2271_t;wire n2272;wire n2272_t;wire n2273;wire n2273_t;wire n2274;wire n2274_t;wire n2275;wire n2275_t;wire n2276;wire n2276_t;wire n2277;wire n2277_t;wire n2278;wire n2278_t;wire n2279;wire n2279_t;wire n2280;wire n2280_t;wire n2281;wire n2281_t;wire n2282;wire n2282_t;wire n2283;wire n2283_t;wire n2284;wire n2284_t;wire n2285;wire n2285_t;wire n2286;wire n2286_t;wire n2287;wire n2287_t;wire n2288;wire n2288_t;wire n2289;wire n2289_t;wire n2290;wire n2290_t;wire n2291;wire n2291_t;wire n2292;wire n2292_t;wire n2293;wire n2293_t;wire n2294;wire n2294_t;wire n2295;wire n2295_t;wire n2296;wire n2296_t;wire n2297;wire n2297_t;wire n2298;wire n2298_t;wire n2299;wire n2299_t;wire n2300;wire n2300_t;wire n2301;wire n2301_t;wire n2302;wire n2302_t;wire n2303;wire n2303_t;wire n2304;wire n2304_t;wire n2307;wire n2307_t;wire n2308;wire n2308_t;wire n2309;wire n2309_t;wire n2310;wire n2310_t;wire n2311;wire n2311_t;wire n2312;wire n2312_t;wire n2313;wire n2313_t;wire n2314;wire n2314_t;wire n2315;wire n2315_t;wire n2316;wire n2316_t;wire n2317;wire n2317_t;wire n2318;wire n2318_t;wire n2319;wire n2319_t;wire n2320;wire n2320_t;wire n2321;wire n2321_t;wire n2322;wire n2322_t;wire n2323;wire n2323_t;wire n2324;wire n2324_t;wire n2325;wire n2325_t;wire n2326;wire n2326_t;wire n2327;wire n2327_t;wire n2328;wire n2328_t;wire n2329;wire n2329_t;wire n2330;wire n2330_t;wire n2331;wire n2331_t;wire n2332;wire n2332_t;wire n2333;wire n2333_t;wire n2334;wire n2334_t;wire n2335;wire n2335_t;wire n2336;wire n2336_t;wire n2337;wire n2337_t;wire n2338;wire n2338_t;wire n2339;wire n2339_t;wire n2340;wire n2340_t;wire n2341;wire n2341_t;wire n2342;wire n2342_t;wire n2343;wire n2343_t;wire n2344;wire n2344_t;wire n2345;wire n2345_t;wire n2346;wire n2346_t;wire n2347;wire n2347_t;wire n2348;wire n2348_t;wire n2349;wire n2349_t;wire n2350;wire n2350_t;wire n2351;wire n2351_t;wire n2352;wire n2352_t;wire n2353;wire n2353_t;wire n2354;wire n2354_t;wire n2355;wire n2355_t;wire n2356;wire n2356_t;wire n2357;wire n2357_t;wire n2358;wire n2358_t;wire n2359;wire n2359_t;wire n2360;wire n2360_t;wire n2361;wire n2361_t;wire n2362;wire n2362_t;wire n2363;wire n2363_t;wire n2364;wire n2364_t;wire n2365;wire n2365_t;wire n2366;wire n2366_t;wire n2367;wire n2367_t;wire n2368;wire n2368_t;wire n2369;wire n2369_t;wire n2370;wire n2370_t;wire n2371;wire n2371_t;wire n2372;wire n2372_t;wire n2373;wire n2373_t;wire n2374;wire n2374_t;wire n2375;wire n2375_t;wire n2376;wire n2376_t;wire n2377;wire n2377_t;wire n2378;wire n2378_t;wire n2379;wire n2379_t;wire n2380;wire n2380_t;wire n2381;wire n2381_t;wire n2382;wire n2382_t;wire n2383;wire n2383_t;wire n2384;wire n2384_t;wire n2385;wire n2385_t;wire n2386;wire n2386_t;wire n2387;wire n2387_t;wire n2388;wire n2388_t;wire n2389;wire n2389_t;wire n2390;wire n2390_t;wire n2391;wire n2391_t;wire n2392;wire n2392_t;wire n2393;wire n2393_t;wire n2394;wire n2394_t;wire n2395;wire n2395_t;wire n2396;wire n2396_t;wire n2397;wire n2397_t;wire n2398;wire n2398_t;wire n2399;wire n2399_t;wire n2400;wire n2400_t;wire n2401;wire n2401_t;wire n2402;wire n2402_t;wire n2403;wire n2403_t;wire n2404;wire n2404_t;wire n2405;wire n2405_t;wire n2406;wire n2406_t;wire n2407;wire n2407_t;wire n2408;wire n2408_t;wire n2409;wire n2409_t;wire n2410;wire n2410_t;wire n2411;wire n2411_t;wire n2412;wire n2412_t;wire n2413;wire n2413_t;wire n2414;wire n2414_t;wire n2415;wire n2415_t;wire n2416;wire n2416_t;wire n2417;wire n2417_t;wire n2418;wire n2418_t;wire n2419;wire n2419_t;wire n2420;wire n2420_t;wire n2421;wire n2421_t;wire n2422;wire n2422_t;wire n2423;wire n2423_t;wire n2424;wire n2424_t;wire n2425;wire n2425_t;wire n2426;wire n2426_t;wire n2427;wire n2427_t;wire n2428;wire n2428_t;wire n2429;wire n2429_t;wire n2430;wire n2430_t;wire n2431;wire n2431_t;wire n2432;wire n2432_t;wire n2433;wire n2433_t;wire n2434;wire n2434_t;wire n2435;wire n2435_t;wire n2436;wire n2436_t;wire n2437;wire n2437_t;wire n2438;wire n2438_t;wire n2439;wire n2439_t;wire n2440;wire n2440_t;wire n2441;wire n2441_t;wire n2442;wire n2442_t;wire n2443;wire n2443_t;wire n2444;wire n2444_t;wire n2445;wire n2445_t;wire n2446;wire n2446_t;wire n2447;wire n2447_t;wire n2448;wire n2448_t;wire n2449;wire n2449_t;wire n2450;wire n2450_t;wire n2451;wire n2451_t;wire n2452;wire n2452_t;wire n2453;wire n2453_t;wire n2454;wire n2454_t;wire n2455;wire n2455_t;wire n2456;wire n2456_t;wire n2457;wire n2457_t;wire n2458;wire n2458_t;wire n2459;wire n2459_t;wire n2460;wire n2460_t;wire n2461;wire n2461_t;wire n2462;wire n2462_t;wire n2463;wire n2463_t;wire n2464;wire n2464_t;wire n2465;wire n2465_t;wire n2466;wire n2466_t;wire n2467;wire n2467_t;wire n2468;wire n2468_t;wire n2469;wire n2469_t;wire n2470;wire n2470_t;wire n2471;wire n2471_t;wire n2472;wire n2472_t;wire n2473;wire n2473_t;wire n2474;wire n2474_t;wire n2475;wire n2475_t;wire n2476;wire n2476_t;wire n2477;wire n2477_t;wire n2478;wire n2478_t;wire n2479;wire n2479_t;wire n2480;wire n2480_t;wire n2481;wire n2481_t;wire n2482;wire n2482_t;wire n2483;wire n2483_t;wire n2484;wire n2484_t;wire n2485;wire n2485_t;wire n2486;wire n2486_t;wire n2487;wire n2487_t;wire n2488;wire n2488_t;wire n2489;wire n2489_t;wire n2490;wire n2490_t;wire n2491;wire n2491_t;wire n2492;wire n2492_t;wire n2493;wire n2493_t;wire n2494;wire n2494_t;wire n2495;wire n2495_t;wire n2496;wire n2496_t;wire n2497;wire n2497_t;wire n2498;wire n2498_t;wire n2499;wire n2499_t;wire n2500;wire n2500_t;wire n2501;wire n2501_t;wire n2502;wire n2502_t;wire n2503;wire n2503_t;wire n2504;wire n2504_t;wire n2505;wire n2505_t;wire n2506;wire n2506_t;wire n2507;wire n2507_t;wire n2508;wire n2508_t;wire n2509;wire n2509_t;wire n2510;wire n2510_t;wire n2511;wire n2511_t;wire n2512;wire n2512_t;wire n2513;wire n2513_t;wire n2514;wire n2514_t;wire n2515;wire n2515_t;wire n2516;wire n2516_t;wire n2517;wire n2517_t;wire n2518;wire n2518_t;wire n2519;wire n2519_t;wire n2520;wire n2520_t;wire n2521;wire n2521_t;wire n2522;wire n2522_t;wire n2523;wire n2523_t;wire n2524;wire n2524_t;wire n2525;wire n2525_t;wire n2526;wire n2526_t;wire n2527;wire n2527_t;wire n2528;wire n2528_t;wire n2529;wire n2529_t;wire n2530;wire n2530_t;wire n2531;wire n2531_t;wire n2532;wire n2532_t;wire n2533;wire n2533_t;wire n2534;wire n2534_t;wire n2535;wire n2535_t;wire n2536;wire n2536_t;wire n2537;wire n2537_t;wire n2538;wire n2538_t;wire n2539;wire n2539_t;wire n2540;wire n2540_t;wire n2541;wire n2541_t;wire n2542;wire n2542_t;wire n2543;wire n2543_t;wire n2544;wire n2544_t;wire n2545;wire n2545_t;wire n2546;wire n2546_t;wire n2547;wire n2547_t;wire n2548;wire n2548_t;wire n2549;wire n2549_t;wire n2550;wire n2550_t;wire n2551;wire n2551_t;wire n2552;wire n2552_t;wire n2553;wire n2553_t;wire n2554;wire n2554_t;wire n2555;wire n2555_t;wire n2556;wire n2556_t;wire n2557;wire n2557_t;wire n2558;wire n2558_t;wire n2559;wire n2559_t;wire n2560;wire n2560_t;wire n2561;wire n2561_t;wire n2562;wire n2562_t;wire n2563;wire n2563_t;wire n2564;wire n2564_t;wire n2565;wire n2565_t;wire n2566;wire n2566_t;wire n2567;wire n2567_t;wire n2568;wire n2568_t;wire n2569;wire n2569_t;wire n2570;wire n2570_t;wire n2571;wire n2571_t;wire n2572;wire n2572_t;wire n2573;wire n2573_t;wire n2574;wire n2574_t;wire n2575;wire n2575_t;wire n2576;wire n2576_t;wire n2577;wire n2577_t;wire n2578;wire n2578_t;wire n2579;wire n2579_t;wire n2580;wire n2580_t;wire n2581;wire n2581_t;wire n2582;wire n2582_t;wire n2583;wire n2583_t;wire n2584;wire n2584_t;wire n2585;wire n2585_t;wire n2586;wire n2586_t;wire n2587;wire n2587_t;wire n2588;wire n2588_t;wire n2589;wire n2589_t;wire n2590;wire n2590_t;wire n2591;wire n2591_t;wire n2592;wire n2592_t;wire n2593;wire n2593_t;wire n2594;wire n2594_t;wire n2595;wire n2595_t;wire n2596;wire n2596_t;wire n2597;wire n2597_t;wire n2598;wire n2598_t;wire n2599;wire n2599_t;wire n2600;wire n2600_t;wire n2601;wire n2601_t;wire n2602;wire n2602_t;wire n2603;wire n2603_t;wire n2604;wire n2604_t;wire n2605;wire n2605_t;wire n2606;wire n2606_t;wire n2607;wire n2607_t;wire n2608;wire n2608_t;wire n2609;wire n2609_t;wire n2610;wire n2610_t;wire n2611;wire n2611_t;wire n2612;wire n2612_t;wire n2613;wire n2613_t;wire n2614;wire n2614_t;wire n2615;wire n2615_t;wire n2616;wire n2616_t;wire n2617;wire n2617_t;wire n2618;wire n2618_t;wire n2619;wire n2619_t;wire n2620;wire n2620_t;wire n2621;wire n2621_t;wire n2622;wire n2622_t;wire n2623;wire n2623_t;wire n2624;wire n2624_t;wire n2625;wire n2625_t;wire n2626;wire n2626_t;wire n2627;wire n2627_t;wire n2628;wire n2628_t;wire n2629;wire n2629_t;wire n2630;wire n2630_t;wire n2631;wire n2631_t;wire n2632;wire n2632_t;wire n2633;wire n2633_t;wire n2634;wire n2634_t;wire n2635;wire n2635_t;wire n2636;wire n2636_t;wire n2637;wire n2637_t;wire n2638;wire n2638_t;wire n2639;wire n2639_t;wire n2640;wire n2640_t;wire n2641;wire n2641_t;wire n2642;wire n2642_t;wire n2643;wire n2643_t;wire n2644;wire n2644_t;wire n2645;wire n2645_t;wire n2646;wire n2646_t;wire n2647;wire n2647_t;wire n2648;wire n2648_t;wire n2649;wire n2649_t;wire n2650;wire n2650_t;wire n2651;wire n2651_t;wire n2652;wire n2652_t;wire n2653;wire n2653_t;wire n2654;wire n2654_t;wire n2655;wire n2655_t;wire n2656;wire n2656_t;wire n2657;wire n2657_t;wire n2658;wire n2658_t;wire n2659;wire n2659_t;wire n2660;wire n2660_t;wire n2661;wire n2661_t;wire n2662;wire n2662_t;wire n2663;wire n2663_t;wire n2664;wire n2664_t;wire n2665;wire n2665_t;wire n2666;wire n2666_t;wire n2667;wire n2667_t;wire n2668;wire n2668_t;wire n2669;wire n2669_t;wire n2670;wire n2670_t;wire n2671;wire n2671_t;wire n2672;wire n2672_t;wire n2673;wire n2673_t;wire n2674;wire n2674_t;wire n2675;wire n2675_t;wire n2676;wire n2676_t;wire n2677;wire n2677_t;wire n2678;wire n2678_t;wire n2679;wire n2679_t;wire n2680;wire n2680_t;wire n2681;wire n2681_t;wire n2682;wire n2682_t;wire n2683;wire n2683_t;wire n2684;wire n2684_t;wire n2685;wire n2685_t;wire n2686;wire n2686_t;wire n2687;wire n2687_t;wire n2688;wire n2688_t;wire n2689;wire n2689_t;wire n2690;wire n2690_t;wire n2691;wire n2691_t;wire n2692;wire n2692_t;wire n2693;wire n2693_t;wire n2694;wire n2694_t;wire n2695;wire n2695_t;wire n2696;wire n2696_t;wire n2697;wire n2697_t;wire n2698;wire n2698_t;wire n2699;wire n2699_t;wire n2700;wire n2700_t;wire n2701;wire n2701_t;wire n2702;wire n2702_t;wire n2703;wire n2703_t;wire n2704;wire n2704_t;wire n2705;wire n2705_t;wire n2706;wire n2706_t;wire n2707;wire n2707_t;wire n2708;wire n2708_t;wire n2709;wire n2709_t;wire n2710;wire n2710_t;wire n2711;wire n2711_t;wire n2712;wire n2712_t;wire n2713;wire n2713_t;wire n2714;wire n2714_t;wire n2715;wire n2715_t;wire n2716;wire n2716_t;wire n2717;wire n2717_t;wire n2718;wire n2718_t;wire n2719;wire n2719_t;wire n2720;wire n2720_t;wire n2721;wire n2721_t;wire n2722;wire n2722_t;wire n2723;wire n2723_t;wire n2724;wire n2724_t;wire n2725;wire n2725_t;wire n2726;wire n2726_t;wire n2727;wire n2727_t;wire n2728;wire n2728_t;wire n2729;wire n2729_t;wire n2730;wire n2730_t;wire n2731;wire n2731_t;wire n2732;wire n2732_t;wire n2733;wire n2733_t;wire n2734;wire n2734_t;wire n2735;wire n2735_t;wire n2736;wire n2736_t;wire n2737;wire n2737_t;wire n2738;wire n2738_t;wire n2739;wire n2739_t;wire n2740;wire n2740_t;wire n2741;wire n2741_t;wire n2742;wire n2742_t;wire n2743;wire n2743_t;wire n2744;wire n2744_t;wire n2745;wire n2745_t;wire n2746;wire n2746_t;wire n2747;wire n2747_t;wire n2748;wire n2748_t;wire n2749;wire n2749_t;wire n2750;wire n2750_t;wire n2751;wire n2751_t;wire n2752;wire n2752_t;wire n2753;wire n2753_t;wire n2754;wire n2754_t;wire n2755;wire n2755_t;wire n2756;wire n2756_t;wire n2757;wire n2757_t;wire n2758;wire n2758_t;wire n2759;wire n2759_t;wire n2760;wire n2760_t;wire n2761;wire n2761_t;wire n2762;wire n2762_t;wire n2763;wire n2763_t;wire n2764;wire n2764_t;wire n2765;wire n2765_t;wire n2766;wire n2766_t;wire n2767;wire n2767_t;wire n2768;wire n2768_t;wire n2769;wire n2769_t;wire n2770;wire n2770_t;wire n2771;wire n2771_t;wire n2772;wire n2772_t;wire n2773;wire n2773_t;wire n2774;wire n2774_t;wire n2775;wire n2775_t;wire n2776;wire n2776_t;wire n2777;wire n2777_t;wire n2778;wire n2778_t;wire n2779;wire n2779_t;wire n2780;wire n2780_t;wire n2781;wire n2781_t;wire n2782;wire n2782_t;wire n2783;wire n2783_t;wire n2784;wire n2784_t;wire n2785;wire n2785_t;wire n2786;wire n2786_t;wire n2787;wire n2787_t;wire n2788;wire n2788_t;wire n2789;wire n2789_t;wire n2790;wire n2790_t;wire n2791;wire n2791_t;wire n2792;wire n2792_t;wire n2793;wire n2793_t;wire n2794;wire n2794_t;wire n2795;wire n2795_t;wire n2796;wire n2796_t;wire n2797;wire n2797_t;wire n2798;wire n2798_t;wire n2799;wire n2799_t;wire n2800;wire n2800_t;wire n2801;wire n2801_t;wire n2802;wire n2802_t;wire n2803;wire n2803_t;wire n2804;wire n2804_t;wire n2805;wire n2805_t;wire n2806;wire n2806_t;wire n2807;wire n2807_t;wire n2808;wire n2808_t;wire n2809;wire n2809_t;wire n2810;wire n2810_t;wire n2811;wire n2811_t;wire n2812;wire n2812_t;wire n2813;wire n2813_t;wire n2814;wire n2814_t;wire n2815;wire n2815_t;wire n2816;wire n2816_t;wire n2817;wire n2817_t;wire n2818;wire n2818_t;wire n2819;wire n2819_t;wire n2820;wire n2820_t;wire n2821;wire n2821_t;wire n2822;wire n2822_t;wire n2823;wire n2823_t;wire n2824;wire n2824_t;wire n2825;wire n2825_t;wire n2826;wire n2826_t;wire n2827;wire n2827_t;wire n2828;wire n2828_t;wire n2829;wire n2829_t;wire n2830;wire n2830_t;wire n2831;wire n2831_t;wire n2832;wire n2832_t;wire n2833;wire n2833_t;wire n2834;wire n2834_t;wire n2835;wire n2835_t;wire n2836;wire n2836_t;wire n2837;wire n2837_t;wire n2838;wire n2838_t;wire n2839;wire n2839_t;wire n2840;wire n2840_t;wire n2841;wire n2841_t;wire n2842;wire n2842_t;wire n2843;wire n2843_t;wire n2844;wire n2844_t;wire n2845;wire n2845_t;wire n2846;wire n2846_t;wire n2847;wire n2847_t;wire n2848;wire n2848_t;wire n2849;wire n2849_t;wire n2850;wire n2850_t;wire n2851;wire n2851_t;wire n2852;wire n2852_t;wire n2853;wire n2853_t;wire n2854;wire n2854_t;wire n2855;wire n2855_t;wire n2856;wire n2856_t;wire n2857;wire n2857_t;wire n2858;wire n2858_t;wire n2859;wire n2859_t;wire n2860;wire n2860_t;wire n2861;wire n2861_t;wire n2862;wire n2862_t;wire n2863;wire n2863_t;wire n2864;wire n2864_t;wire n2865;wire n2865_t;wire n2866;wire n2866_t;wire n2867;wire n2867_t;wire n2868;wire n2868_t;wire n2869;wire n2869_t;wire n2870;wire n2870_t;wire n2871;wire n2871_t;wire n2872;wire n2872_t;wire n2873;wire n2873_t;wire n2874;wire n2874_t;wire n2875;wire n2875_t;wire n2876;wire n2876_t;wire n2877;wire n2877_t;wire n2878;wire n2878_t;wire n2879;wire n2879_t;wire n2880;wire n2880_t;wire n2881;wire n2881_t;wire n2882;wire n2882_t;wire n2883;wire n2883_t;wire n2884;wire n2884_t;wire n2885;wire n2885_t;wire n2886;wire n2886_t;wire n2887;wire n2887_t;wire n2888;wire n2888_t;wire n2889;wire n2889_t;wire n2890;wire n2890_t;wire n2891;wire n2891_t;wire n2892;wire n2892_t;wire n2893;wire n2893_t;wire n2894;wire n2894_t;wire n2895;wire n2895_t;wire n2896;wire n2896_t;wire n2897;wire n2897_t;wire n2898;wire n2898_t;wire n2899;wire n2899_t;wire n2900;wire n2900_t;wire n2901;wire n2901_t;wire n2902;wire n2902_t;wire n2903;wire n2903_t;wire n2904;wire n2904_t;wire n2905;wire n2905_t;wire n2906;wire n2906_t;wire n2907;wire n2907_t;wire n2908;wire n2908_t;wire n2909;wire n2909_t;wire n2910;wire n2910_t;wire n2911;wire n2911_t;wire n2912;wire n2912_t;wire n2913;wire n2913_t;wire n2914;wire n2914_t;wire n2915;wire n2915_t;wire n2916;wire n2916_t;wire n2917;wire n2917_t;wire n2918;wire n2918_t;wire n2919;wire n2919_t;wire n2920;wire n2920_t;wire n2921;wire n2921_t;wire n2922;wire n2922_t;wire n2923;wire n2923_t;wire n2924;wire n2924_t;wire n2925;wire n2925_t;wire n2926;wire n2926_t;wire n2927;wire n2927_t;wire n2928;wire n2928_t;wire n2929;wire n2929_t;wire n2930;wire n2930_t;wire n2931;wire n2931_t;wire n2932;wire n2932_t;wire n2933;wire n2933_t;wire n2934;wire n2934_t;wire n2935;wire n2935_t;wire n2936;wire n2936_t;wire n2937;wire n2937_t;wire n2938;wire n2938_t;wire n2939;wire n2939_t;wire n2940;wire n2940_t;wire n2941;wire n2941_t;wire n2942;wire n2942_t;wire n2943;wire n2943_t;wire n2944;wire n2944_t;wire n2945;wire n2945_t;wire n2946;wire n2946_t;wire n2947;wire n2947_t;wire n2948;wire n2948_t;wire n2949;wire n2949_t;wire n2950;wire n2950_t;wire n2951;wire n2951_t;wire n2952;wire n2952_t;wire n2953;wire n2953_t;wire n2954;wire n2954_t;wire n2955;wire n2955_t;wire n2956;wire n2956_t;wire n2957;wire n2957_t;wire n2958;wire n2958_t;wire n2959;wire n2959_t;wire n2960;wire n2960_t;wire n2961;wire n2961_t;wire n2962;wire n2962_t;wire n2963;wire n2963_t;wire n2964;wire n2964_t;wire n2965;wire n2965_t;wire n2966;wire n2966_t;wire n2967;wire n2967_t;wire n2968;wire n2968_t;wire n2969;wire n2969_t;wire n2970;wire n2970_t;wire n2971;wire n2971_t;wire n2972;wire n2972_t;wire n2973;wire n2973_t;wire n2974;wire n2974_t;wire n2975;wire n2975_t;wire n2976;wire n2976_t;wire n2977;wire n2977_t;wire n2978;wire n2978_t;wire n2979;wire n2979_t;wire n2980;wire n2980_t;wire n2981;wire n2981_t;wire n2982;wire n2982_t;wire n2983;wire n2983_t;wire n2984;wire n2984_t;wire n2985;wire n2985_t;wire n2986;wire n2986_t;wire n2987;wire n2987_t;wire n2988;wire n2988_t;wire n2989;wire n2989_t;wire n2990;wire n2990_t;wire n2991;wire n2991_t;wire n2992;wire n2992_t;wire n2993;wire n2993_t;wire n2994;wire n2994_t;wire n2995;wire n2995_t;wire n2996;wire n2996_t;wire n2997;wire n2997_t;wire n2998;wire n2998_t;wire n2999;wire n2999_t;wire n3000;wire n3000_t;wire n3001;wire n3001_t;wire n3002;wire n3002_t;wire n3003;wire n3003_t;wire n3004;wire n3004_t;wire n3005;wire n3005_t;wire n3006;wire n3006_t;wire n3007;wire n3007_t;wire n3008;wire n3008_t;wire n3009;wire n3009_t;wire n3010;wire n3010_t;wire n3011;wire n3011_t;wire n3012;wire n3012_t;wire n3013;wire n3013_t;wire n3014;wire n3014_t;wire n3015;wire n3015_t;wire n3016;wire n3016_t;wire n3017;wire n3017_t;wire n3018;wire n3018_t;wire n3019;wire n3019_t;wire n3020;wire n3020_t;wire n3021;wire n3021_t;wire n3022;wire n3022_t;wire n3023;wire n3023_t;wire n3024;wire n3024_t;wire n3025;wire n3025_t;wire n3026;wire n3026_t;wire n3027;wire n3027_t;wire n3028;wire n3028_t;wire n3029;wire n3029_t;wire n3030;wire n3030_t;wire n3031;wire n3031_t;wire n3032;wire n3032_t;wire n3033;wire n3033_t;wire n3034;wire n3034_t;wire n3035;wire n3035_t;wire n3036;wire n3036_t;wire n3037;wire n3037_t;wire n3038;wire n3038_t;wire n3039;wire n3039_t;wire n3040;wire n3040_t;wire n3041;wire n3041_t;wire n3042;wire n3042_t;wire n3043;wire n3043_t;wire n3044;wire n3044_t;wire n3045;wire n3045_t;wire n3046;wire n3046_t;wire n3047;wire n3047_t;wire n3048;wire n3048_t;wire n3049;wire n3049_t;wire n3050;wire n3050_t;wire n3051;wire n3051_t;wire n3052;wire n3052_t;wire n3053;wire n3053_t;wire n3054;wire n3054_t;wire n3055;wire n3055_t;wire n3056;wire n3056_t;wire n3057;wire n3057_t;wire n3058;wire n3058_t;wire n3059;wire n3059_t;wire n3060;wire n3060_t;wire n3061;wire n3061_t;wire n3062;wire n3062_t;wire n3063;wire n3063_t;wire n3064;wire n3064_t;wire n3065;wire n3065_t;wire n3066;wire n3066_t;wire n3067;wire n3067_t;wire n3068;wire n3068_t;wire n3069;wire n3069_t;wire n3070;wire n3070_t;wire n3071;wire n3071_t;wire n3072;wire n3072_t;wire n3073;wire n3073_t;wire n3074;wire n3074_t;wire n3075;wire n3075_t;wire n3076;wire n3076_t;wire n3077;wire n3077_t;wire n3078;wire n3078_t;wire n3079;wire n3079_t;wire n3080;wire n3080_t;wire n3081;wire n3081_t;wire n3082;wire n3082_t;wire n3083;wire n3083_t;wire n3084;wire n3084_t;wire n3085;wire n3085_t;wire n3086;wire n3086_t;wire n3087;wire n3087_t;wire n3088;wire n3088_t;wire n3089;wire n3089_t;wire n3090;wire n3090_t;wire n3091;wire n3091_t;wire n3092;wire n3092_t;wire n3093;wire n3093_t;wire n3094;wire n3094_t;wire n3095;wire n3095_t;wire n3096;wire n3096_t;wire n3097;wire n3097_t;wire n3098;wire n3098_t;wire n3099;wire n3099_t;wire n3100;wire n3100_t;wire n3101;wire n3101_t;wire n3102;wire n3102_t;wire n3103;wire n3103_t;wire n3104;wire n3104_t;wire n3105;wire n3105_t;wire n3106;wire n3106_t;wire n3107;wire n3107_t;wire n3108;wire n3108_t;wire n3109;wire n3109_t;wire n3110;wire n3110_t;wire n3111;wire n3111_t;wire n3112;wire n3112_t;wire n3113;wire n3113_t;wire n3114;wire n3114_t;wire n3115;wire n3115_t;wire n3116;wire n3116_t;wire n3117;wire n3117_t;wire n3118;wire n3118_t;wire n3119;wire n3119_t;wire n3120;wire n3120_t;wire n3121;wire n3121_t;wire n3122;wire n3122_t;wire n3123;wire n3123_t;wire n3124;wire n3124_t;wire n3125;wire n3125_t;wire n3126;wire n3126_t;wire n3127;wire n3127_t;wire n3128;wire n3128_t;wire n3129;wire n3129_t;wire n3130;wire n3130_t;wire n3131;wire n3131_t;wire n3132;wire n3132_t;wire n3133;wire n3133_t;wire n3134;wire n3134_t;wire n3135;wire n3135_t;wire n3136;wire n3136_t;wire n3137;wire n3137_t;wire n3138;wire n3138_t;wire n3139;wire n3139_t;wire n3140;wire n3140_t;wire n3141;wire n3141_t;wire n3142;wire n3142_t;wire n3143;wire n3143_t;wire n3144;wire n3144_t;wire n3145;wire n3145_t;wire n3146;wire n3146_t;wire n3147;wire n3147_t;wire n3148;wire n3148_t;wire n3149;wire n3149_t;wire n3150;wire n3150_t;wire n3151;wire n3151_t;wire n3152;wire n3152_t;wire n3153;wire n3153_t;wire n3154;wire n3154_t;wire n3155;wire n3155_t;wire n3156;wire n3156_t;wire n3157;wire n3157_t;wire n3158;wire n3158_t;wire n3159;wire n3159_t;wire n3160;wire n3160_t;wire n3161;wire n3161_t;wire n3162;wire n3162_t;wire n3163;wire n3163_t;wire n3164;wire n3164_t;wire n3165;wire n3165_t;wire n3166;wire n3166_t;wire n3167;wire n3167_t;wire n3168;wire n3168_t;wire n3169;wire n3169_t;wire n3170;wire n3170_t;wire n3171;wire n3171_t;wire n3172;wire n3172_t;wire n3173;wire n3173_t;wire n3174;wire n3174_t;wire n3175;wire n3175_t;wire n3176;wire n3176_t;wire n3177;wire n3177_t;wire n3178;wire n3178_t;wire n3179;wire n3179_t;wire n3180;wire n3180_t;wire n3181;wire n3181_t;wire n3182;wire n3182_t;wire n3183;wire n3183_t;wire n3184;wire n3184_t;wire n3185;wire n3185_t;wire n3186;wire n3186_t;wire n3187;wire n3187_t;wire n3188;wire n3188_t;wire n3189;wire n3189_t;wire n3190;wire n3190_t;wire n3191;wire n3191_t;wire n3192;wire n3192_t;wire n3193;wire n3193_t;wire n3194;wire n3194_t;wire n3195;wire n3195_t;wire n3196;wire n3196_t;wire n3197;wire n3197_t;wire n3198;wire n3198_t;wire n3199;wire n3199_t;wire n3200;wire n3200_t;wire n3201;wire n3201_t;wire n3202;wire n3202_t;wire n3203;wire n3203_t;wire n3204;wire n3204_t;wire n3333;wire n3333_t;wire n3334;wire n3334_t;wire n3335;wire n3335_t;wire n3336;wire n3336_t;wire n3337;wire n3337_t;wire n3338;wire n3338_t;wire n3339;wire n3339_t;wire n3340;wire n3340_t;wire n3341;wire n3341_t;wire n3342;wire n3342_t;wire n3343;wire n3343_t;wire n3344;wire n3344_t;wire n3345;wire n3345_t;wire n3346;wire n3346_t;wire n3347;wire n3347_t;wire n3348;wire n3348_t;wire n3349;wire n3349_t;wire n3350;wire n3350_t;wire n3351;wire n3351_t;wire n3352;wire n3352_t;wire n3353;wire n3353_t;wire n3354;wire n3354_t;wire n3355;wire n3355_t;wire n3356;wire n3356_t;wire n3357;wire n3357_t;wire n3358;wire n3358_t;wire n3359;wire n3359_t;wire n3360;wire n3360_t;wire n3361;wire n3361_t;wire n3362;wire n3362_t;wire n3363;wire n3363_t;wire n3364;wire n3364_t;wire n3365;wire n3365_t;wire n3366;wire n3366_t;wire n3367;wire n3367_t;wire n3368;wire n3368_t;wire n3369;wire n3369_t;wire n3370;wire n3370_t;wire n3371;wire n3371_t;wire n3372;wire n3372_t;wire n3373;wire n3373_t;wire n3374;wire n3374_t;wire n3375;wire n3375_t;wire n3376;wire n3376_t;wire n3377;wire n3377_t;wire n3378;wire n3378_t;wire n3379;wire n3379_t;wire n3380;wire n3380_t;wire n3381;wire n3381_t;wire n3382;wire n3382_t;wire n3383;wire n3383_t;wire n3384;wire n3384_t;wire n3385;wire n3385_t;wire n3386;wire n3386_t;wire n3387;wire n3387_t;wire n3388;wire n3388_t;wire n3389;wire n3389_t;wire n3390;wire n3390_t;wire n3391;wire n3391_t;wire n3392;wire n3392_t;wire n3393;wire n3393_t;wire n3394;wire n3394_t;wire n3395;wire n3395_t;wire n3396;wire n3396_t;wire n3397;wire n3397_t;wire n3398;wire n3398_t;wire n3399;wire n3399_t;wire n3400;wire n3400_t;wire n3401;wire n3401_t;wire n3402;wire n3402_t;wire n3403;wire n3403_t;wire n3404;wire n3404_t;wire n3405;wire n3405_t;wire n3406;wire n3406_t;wire n3407;wire n3407_t;wire n3408;wire n3408_t;wire n3409;wire n3409_t;wire n3410;wire n3410_t;wire n3411;wire n3411_t;wire n3412;wire n3412_t;wire n3413;wire n3413_t;wire n3414;wire n3414_t;wire n3415;wire n3415_t;wire n3416;wire n3416_t;wire n3417;wire n3417_t;wire n3418;wire n3418_t;wire n3419;wire n3419_t;wire n3420;wire n3420_t;wire n3421;wire n3421_t;wire n3422;wire n3422_t;wire n3423;wire n3423_t;wire n3424;wire n3424_t;wire n3425;wire n3425_t;wire n3426;wire n3426_t;wire n3427;wire n3427_t;wire n3428;wire n3428_t;wire n3429;wire n3429_t;wire n3430;wire n3430_t;wire n3431;wire n3431_t;wire n3432;wire n3432_t;wire n3433;wire n3433_t;wire n3434;wire n3434_t;wire n3435;wire n3435_t;wire n3436;wire n3436_t;wire n3437;wire n3437_t;wire n3438;wire n3438_t;wire n3439;wire n3439_t;wire n3440;wire n3440_t;wire n3441;wire n3441_t;wire n3442;wire n3442_t;wire n3443;wire n3443_t;wire n3444;wire n3444_t;wire n3445;wire n3445_t;wire n3446;wire n3446_t;wire n3447;wire n3447_t;wire n3448;wire n3448_t;wire n3449;wire n3449_t;wire n3450;wire n3450_t;wire n3451;wire n3451_t;wire n3452;wire n3452_t;wire n3453;wire n3453_t;wire n3454;wire n3454_t;wire n3455;wire n3455_t;wire n3456;wire n3456_t;wire n3457;wire n3457_t;wire n3458;wire n3458_t;wire n3459;wire n3459_t;wire n3460;wire n3460_t;wire n3461;wire n3461_t;wire n3462;wire n3462_t;wire n3463;wire n3463_t;wire n3464;wire n3464_t;wire n3465;wire n3465_t;wire n3466;wire n3466_t;wire n3467;wire n3467_t;wire n3468;wire n3468_t;wire n3469;wire n3469_t;wire n3470;wire n3470_t;wire n3471;wire n3471_t;wire n3472;wire n3472_t;wire n3473;wire n3473_t;wire n3474;wire n3474_t;wire n3475;wire n3475_t;wire n3476;wire n3476_t;wire n3477;wire n3477_t;wire n3478;wire n3478_t;wire n3479;wire n3479_t;wire n3480;wire n3480_t;wire n3481;wire n3481_t;wire n3482;wire n3482_t;wire n3483;wire n3483_t;wire n3484;wire n3484_t;wire n3485;wire n3485_t;wire n3486;wire n3486_t;wire n3487;wire n3487_t;wire n3488;wire n3488_t;wire n3489;wire n3489_t;wire n3490;wire n3490_t;wire n3491;wire n3491_t;wire n3492;wire n3492_t;wire n3493;wire n3493_t;wire n3494;wire n3494_t;wire n3495;wire n3495_t;wire n3496;wire n3496_t;wire n3497;wire n3497_t;wire n3498;wire n3498_t;wire n3499;wire n3499_t;wire n3500;wire n3500_t;wire n3501;wire n3501_t;wire n3502;wire n3502_t;wire n3503;wire n3503_t;wire n3504;wire n3504_t;wire n3505;wire n3505_t;wire n3506;wire n3506_t;wire n3507;wire n3507_t;wire n3508;wire n3508_t;wire n3509;wire n3509_t;wire n3510;wire n3510_t;wire n3511;wire n3511_t;wire n3512;wire n3512_t;wire n3513;wire n3513_t;wire n3514;wire n3514_t;wire n3515;wire n3515_t;wire n3516;wire n3516_t;wire n3517;wire n3517_t;wire n3518;wire n3518_t;wire n3519;wire n3519_t;wire n3520;wire n3520_t;wire n3521;wire n3521_t;wire n3522;wire n3522_t;wire n3523;wire n3523_t;wire n3524;wire n3524_t;wire n3525;wire n3525_t;wire n3526;wire n3526_t;wire n3527;wire n3527_t;wire n3528;wire n3528_t;wire n3529;wire n3529_t;wire n3530;wire n3530_t;wire n3531;wire n3531_t;wire n3532;wire n3532_t;wire n3533;wire n3533_t;wire n3534;wire n3534_t;wire n3535;wire n3535_t;wire n3536;wire n3536_t;wire n3537;wire n3537_t;wire n3538;wire n3538_t;wire n3539;wire n3539_t;wire n3540;wire n3540_t;wire n3541;wire n3541_t;wire n3542;wire n3542_t;wire n3543;wire n3543_t;wire n3544;wire n3544_t;wire n3545;wire n3545_t;wire n3546;wire n3546_t;wire n3547;wire n3547_t;wire n3548;wire n3548_t;wire n3549;wire n3549_t;wire n3550;wire n3550_t;wire n3551;wire n3551_t;wire n3552;wire n3552_t;wire n3553;wire n3553_t;wire n3554;wire n3554_t;wire n3555;wire n3555_t;wire n3556;wire n3556_t;wire n3557;wire n3557_t;wire n3558;wire n3558_t;wire n3559;wire n3559_t;wire n3560;wire n3560_t;wire n3561;wire n3561_t;wire n3562;wire n3562_t;wire n3563;wire n3563_t;wire n3564;wire n3564_t;wire n3565;wire n3565_t;wire n3566;wire n3566_t;wire n3567;wire n3567_t;wire n3568;wire n3568_t;wire n3569;wire n3569_t;wire n3570;wire n3570_t;wire n3571;wire n3571_t;wire n3572;wire n3572_t;wire n3573;wire n3573_t;wire n3574;wire n3574_t;wire n3575;wire n3575_t;wire n3576;wire n3576_t;wire n3577;wire n3577_t;wire n3578;wire n3578_t;wire n3579;wire n3579_t;wire n3580;wire n3580_t;wire n3581;wire n3581_t;wire n3582;wire n3582_t;wire n3583;wire n3583_t;wire n3584;wire n3584_t;wire n3585;wire n3585_t;wire n3586;wire n3586_t;wire n3587;wire n3587_t;wire n3588;wire n3588_t;wire n3589;wire n3589_t;wire n3590;wire n3590_t;wire n3591;wire n3591_t;wire n3592;wire n3592_t;wire n3593;wire n3593_t;wire n3594;wire n3594_t;wire n3595;wire n3595_t;wire n3596;wire n3596_t;wire n3597;wire n3597_t;wire n3598;wire n3598_t;wire n3599;wire n3599_t;wire n3600;wire n3600_t;wire n3601;wire n3601_t;wire n3602;wire n3602_t;wire n3603;wire n3603_t;wire n3604;wire n3604_t;wire n3605;wire n3605_t;wire n3606;wire n3606_t;wire n3607;wire n3607_t;wire n3608;wire n3608_t;wire n3609;wire n3609_t;wire n3610;wire n3610_t;wire n3611;wire n3611_t;wire n3612;wire n3612_t;wire n3613;wire n3613_t;wire n3614;wire n3614_t;wire n3615;wire n3615_t;wire n3616;wire n3616_t;wire n3617;wire n3617_t;wire n3618;wire n3618_t;wire n3619;wire n3619_t;wire n3620;wire n3620_t;wire n3621;wire n3621_t;wire n3622;wire n3622_t;wire n3623;wire n3623_t;wire n3624;wire n3624_t;wire n3625;wire n3625_t;wire n3626;wire n3626_t;wire n3627;wire n3627_t;wire n3628;wire n3628_t;wire n3629;wire n3629_t;wire n3630;wire n3630_t;wire n3631;wire n3631_t;wire n3632;wire n3632_t;wire n3633;wire n3633_t;wire n3634;wire n3634_t;wire n3635;wire n3635_t;wire n3636;wire n3636_t;wire n3637;wire n3637_t;wire n3638;wire n3638_t;wire n3639;wire n3639_t;wire n3640;wire n3640_t;wire n3641;wire n3641_t;wire n3642;wire n3642_t;wire n3643;wire n3643_t;wire n3644;wire n3644_t;wire n3645;wire n3645_t;wire n3646;wire n3646_t;wire n3647;wire n3647_t;wire n3648;wire n3648_t;wire n3649;wire n3649_t;wire n3650;wire n3650_t;wire n3651;wire n3651_t;wire n3652;wire n3652_t;wire n3653;wire n3653_t;wire n3654;wire n3654_t;wire n3655;wire n3655_t;wire n3656;wire n3656_t;wire n3657;wire n3657_t;wire n3658;wire n3658_t;wire n3659;wire n3659_t;wire n3660;wire n3660_t;wire n3661;wire n3661_t;wire n3662;wire n3662_t;wire n3663;wire n3663_t;wire n3664;wire n3664_t;wire n3665;wire n3665_t;wire n3666;wire n3666_t;wire n3667;wire n3667_t;wire n3668;wire n3668_t;wire n3669;wire n3669_t;wire n3670;wire n3670_t;wire n3671;wire n3671_t;wire n3672;wire n3672_t;wire n3673;wire n3673_t;wire n3674;wire n3674_t;wire n3675;wire n3675_t;wire n3676;wire n3676_t;wire n3677;wire n3677_t;wire n3678;wire n3678_t;wire n3679;wire n3679_t;wire n3680;wire n3680_t;wire n3681;wire n3681_t;wire n3682;wire n3682_t;wire n3683;wire n3683_t;wire n3684;wire n3684_t;wire n3685;wire n3685_t;wire n3686;wire n3686_t;wire n3687;wire n3687_t;wire n3688;wire n3688_t;wire n3689;wire n3689_t;wire n3690;wire n3690_t;wire n3691;wire n3691_t;wire n3692;wire n3692_t;wire n3693;wire n3693_t;wire n3694;wire n3694_t;wire n3695;wire n3695_t;wire n3696;wire n3696_t;wire n3697;wire n3697_t;wire n3698;wire n3698_t;wire n3699;wire n3699_t;wire n3700;wire n3700_t;wire n3701;wire n3701_t;wire n3702;wire n3702_t;wire n3703;wire n3703_t;wire n3704;wire n3704_t;wire n3705;wire n3705_t;wire n3706;wire n3706_t;wire n3707;wire n3707_t;wire n3708;wire n3708_t;wire n3709;wire n3709_t;wire n3710;wire n3710_t;wire n3711;wire n3711_t;wire n3712;wire n3712_t;wire n3713;wire n3713_t;wire n3714;wire n3714_t;wire n3715;wire n3715_t;wire n3716;wire n3716_t;wire n3717;wire n3717_t;wire n3718;wire n3718_t;wire n3719;wire n3719_t;wire n3720;wire n3720_t;wire n3721;wire n3721_t;wire n3722;wire n3722_t;wire n3723;wire n3723_t;wire n3724;wire n3724_t;wire n3725;wire n3725_t;wire n3726;wire n3726_t;wire n3727;wire n3727_t;wire n3728;wire n3728_t;wire n3729;wire n3729_t;wire n3730;wire n3730_t;wire n3731;wire n3731_t;wire n3732;wire n3732_t;wire n3733;wire n3733_t;wire n3734;wire n3734_t;wire n3735;wire n3735_t;wire n3736;wire n3736_t;wire n3737;wire n3737_t;wire n3738;wire n3738_t;wire n3739;wire n3739_t;wire n3740;wire n3740_t;wire n3741;wire n3741_t;wire n3742;wire n3742_t;wire n3743;wire n3743_t;wire n3744;wire n3744_t;wire n3745;wire n3745_t;wire n3746;wire n3746_t;wire n3747;wire n3747_t;wire n3748;wire n3748_t;wire n3749;wire n3749_t;wire n3750;wire n3750_t;wire n3751;wire n3751_t;wire n3752;wire n3752_t;wire n3753;wire n3753_t;wire n3754;wire n3754_t;wire n3755;wire n3755_t;wire n3756;wire n3756_t;wire n3757;wire n3757_t;wire n3758;wire n3758_t;wire n3759;wire n3759_t;wire n3760;wire n3760_t;wire n3761;wire n3761_t;wire n3762;wire n3762_t;wire n3763;wire n3763_t;wire n3764;wire n3764_t;wire n3765;wire n3765_t;wire n3766;wire n3766_t;wire n3767;wire n3767_t;wire n3768;wire n3768_t;wire n3769;wire n3769_t;wire n3770;wire n3770_t;wire n3771;wire n3771_t;wire n3772;wire n3772_t;wire n3773;wire n3773_t;wire n3774;wire n3774_t;wire n3775;wire n3775_t;wire n3776;wire n3776_t;wire n3777;wire n3777_t;wire n3778;wire n3778_t;wire n3779;wire n3779_t;wire n3780;wire n3780_t;wire n3781;wire n3781_t;wire n3782;wire n3782_t;wire n3783;wire n3783_t;wire n3784;wire n3784_t;wire n3785;wire n3785_t;wire n3786;wire n3786_t;wire n3787;wire n3787_t;wire n3788;wire n3788_t;wire n3789;wire n3789_t;wire n3790;wire n3790_t;wire n3791;wire n3791_t;wire n3792;wire n3792_t;wire n3793;wire n3793_t;wire n3794;wire n3794_t;wire n3795;wire n3795_t;wire n3796;wire n3796_t;wire n3797;wire n3797_t;wire n3798;wire n3798_t;wire n3799;wire n3799_t;wire n3800;wire n3800_t;wire n3801;wire n3801_t;wire n3802;wire n3802_t;wire n3803;wire n3803_t;wire n3804;wire n3804_t;wire n3805;wire n3805_t;wire n3806;wire n3806_t;wire n3807;wire n3807_t;wire n3808;wire n3808_t;wire n3809;wire n3809_t;wire n3810;wire n3810_t;wire n3811;wire n3811_t;wire n3812;wire n3812_t;wire n3813;wire n3813_t;wire n3814;wire n3814_t;wire n3815;wire n3815_t;wire n3816;wire n3816_t;wire n3817;wire n3817_t;wire n3818;wire n3818_t;wire n3819;wire n3819_t;wire n3820;wire n3820_t;wire n3821;wire n3821_t;wire n3822;wire n3822_t;wire n3823;wire n3823_t;wire n3824;wire n3824_t;wire n3825;wire n3825_t;wire n3826;wire n3826_t;wire n3827;wire n3827_t;wire n3828;wire n3828_t;wire n3829;wire n3829_t;wire n3830;wire n3830_t;wire n3831;wire n3831_t;wire n3832;wire n3832_t;wire n3833;wire n3833_t;wire n3834;wire n3834_t;wire n3835;wire n3835_t;wire n3836;wire n3836_t;wire n3837;wire n3837_t;wire n3838;wire n3838_t;wire n3839;wire n3839_t;wire n3840;wire n3840_t;wire n3841;wire n3841_t;wire n3842;wire n3842_t;wire n3843;wire n3843_t;wire n3844;wire n3844_t;wire n3845;wire n3845_t;wire n3846;wire n3846_t;wire n3847;wire n3847_t;wire n3848;wire n3848_t;wire n3849;wire n3849_t;wire n3850;wire n3850_t;wire n3851;wire n3851_t;wire n3852;wire n3852_t;wire n3853;wire n3853_t;wire n3854;wire n3854_t;wire n3855;wire n3855_t;wire n3856;wire n3856_t;wire n3857;wire n3857_t;wire n3858;wire n3858_t;wire n3859;wire n3859_t;wire n3860;wire n3860_t;wire n3861;wire n3861_t;wire n3862;wire n3862_t;wire n3863;wire n3863_t;wire n3864;wire n3864_t;wire n3865;wire n3865_t;wire n3866;wire n3866_t;wire n3867;wire n3867_t;wire n3868;wire n3868_t;wire n3869;wire n3869_t;wire n3870;wire n3870_t;wire n3871;wire n3871_t;wire n3872;wire n3872_t;wire n3873;wire n3873_t;wire n3874;wire n3874_t;wire n3875;wire n3875_t;wire n3876;wire n3876_t;wire n3877;wire n3877_t;wire n3878;wire n3878_t;wire n3879;wire n3879_t;wire n3880;wire n3880_t;wire n3881;wire n3881_t;wire n3882;wire n3882_t;wire n3883;wire n3883_t;wire n3884;wire n3884_t;wire n3885;wire n3885_t;wire n3886;wire n3886_t;wire n3887;wire n3887_t;wire n3888;wire n3888_t;wire n3889;wire n3889_t;wire n3890;wire n3890_t;wire n3891;wire n3891_t;wire n3892;wire n3892_t;wire n3893;wire n3893_t;wire n3894;wire n3894_t;wire n3895;wire n3895_t;wire n3896;wire n3896_t;wire n3897;wire n3897_t;wire n3898;wire n3898_t;wire n3899;wire n3899_t;wire n3900;wire n3900_t;wire n3901;wire n3901_t;wire n3902;wire n3902_t;wire n3903;wire n3903_t;wire n3904;wire n3904_t;wire n3905;wire n3905_t;wire n3906;wire n3906_t;wire n3907;wire n3907_t;wire n3908;wire n3908_t;wire n3909;wire n3909_t;wire n3910;wire n3910_t;wire n3911;wire n3911_t;wire n3912;wire n3912_t;wire n3913;wire n3913_t;wire n3914;wire n3914_t;wire n3915;wire n3915_t;wire n3916;wire n3916_t;wire n3917;wire n3917_t;wire n3918;wire n3918_t;wire n3919;wire n3919_t;wire n3920;wire n3920_t;wire n3921;wire n3921_t;wire n3922;wire n3922_t;wire n3923;wire n3923_t;wire n3924;wire n3924_t;wire n3925;wire n3925_t;wire n3926;wire n3926_t;wire n3927;wire n3927_t;wire n3928;wire n3928_t;wire n3929;wire n3929_t;wire n3930;wire n3930_t;wire n3931;wire n3931_t;wire n3932;wire n3932_t;wire n3933;wire n3933_t;wire n3934;wire n3934_t;wire n3935;wire n3935_t;wire n3936;wire n3936_t;wire n3937;wire n3937_t;wire n3938;wire n3938_t;wire n3939;wire n3939_t;wire n3940;wire n3940_t;wire n3941;wire n3941_t;wire n3942;wire n3942_t;wire n3943;wire n3943_t;wire n3944;wire n3944_t;wire n3945;wire n3945_t;wire n3946;wire n3946_t;wire n3947;wire n3947_t;wire n3948;wire n3948_t;wire n3949;wire n3949_t;wire n3950;wire n3950_t;wire n3951;wire n3951_t;wire n3952;wire n3952_t;wire n3953;wire n3953_t;wire n3954;wire n3954_t;wire n3955;wire n3955_t;wire n3956;wire n3956_t;wire n3957;wire n3957_t;wire n3958;wire n3958_t;wire n3959;wire n3959_t;wire n3960;wire n3960_t;wire n3961;wire n3961_t;wire n3962;wire n3962_t;wire n3963;wire n3963_t;wire n3964;wire n3964_t;wire n3965;wire n3965_t;wire n3966;wire n3966_t;wire n3967;wire n3967_t;wire n3968;wire n3968_t;wire n3969;wire n3969_t;wire n3970;wire n3970_t;wire n3971;wire n3971_t;wire n3972;wire n3972_t;wire n3973;wire n3973_t;wire n3974;wire n3974_t;wire n3975;wire n3975_t;wire n3976;wire n3976_t;wire n3977;wire n3977_t;wire n3978;wire n3978_t;wire n3979;wire n3979_t;wire n3980;wire n3980_t;wire n3981;wire n3981_t;wire n3982;wire n3982_t;wire n3983;wire n3983_t;wire n3984;wire n3984_t;wire n3985;wire n3985_t;wire n3986;wire n3986_t;wire n3987;wire n3987_t;wire n3988;wire n3988_t;wire n3989;wire n3989_t;wire n3990;wire n3990_t;wire n3991;wire n3991_t;wire n3992;wire n3992_t;wire n3993;wire n3993_t;wire n3994;wire n3994_t;wire n3995;wire n3995_t;wire n3996;wire n3996_t;wire n3997;wire n3997_t;wire n3998;wire n3998_t;wire n3999;wire n3999_t;wire n4000;wire n4000_t;wire n4001;wire n4001_t;wire n4002;wire n4002_t;wire n4003;wire n4003_t;wire n4004;wire n4004_t;wire n4005;wire n4005_t;wire n4006;wire n4006_t;wire n4007;wire n4007_t;wire n4008;wire n4008_t;wire n4009;wire n4009_t;wire n4010;wire n4010_t;wire n4011;wire n4011_t;wire n4012;wire n4012_t;wire n4013;wire n4013_t;wire n4014;wire n4014_t;wire n4015;wire n4015_t;wire n4016;wire n4016_t;wire n4017;wire n4017_t;wire n4018;wire n4018_t;wire n4019;wire n4019_t;wire n4020;wire n4020_t;wire n4021;wire n4021_t;wire n4022;wire n4022_t;wire n4023;wire n4023_t;wire n4024;wire n4024_t;wire n4025;wire n4025_t;wire n4026;wire n4026_t;wire n4027;wire n4027_t;wire n4028;wire n4028_t;wire n4029;wire n4029_t;wire n4030;wire n4030_t;wire n4031;wire n4031_t;wire n4032;wire n4032_t;wire n4033;wire n4033_t;wire n4034;wire n4034_t;wire n4035;wire n4035_t;wire n4036;wire n4036_t;wire n4037;wire n4037_t;wire n4038;wire n4038_t;wire n4039;wire n4039_t;wire n4040;wire n4040_t;wire n4041;wire n4041_t;wire n4042;wire n4042_t;wire n4043;wire n4043_t;wire n4044;wire n4044_t;wire n4045;wire n4045_t;wire n4046;wire n4046_t;wire n4047;wire n4047_t;wire n4048;wire n4048_t;wire n4049;wire n4049_t;wire n4050;wire n4050_t;wire n4051;wire n4051_t;wire n4052;wire n4052_t;wire n4053;wire n4053_t;wire n4054;wire n4054_t;wire n4055;wire n4055_t;wire n4056;wire n4056_t;wire n4057;wire n4057_t;wire n4058;wire n4058_t;wire n4059;wire n4059_t;wire n4060;wire n4060_t;wire n4061;wire n4061_t;wire n4062;wire n4062_t;wire n4063;wire n4063_t;wire n4064;wire n4064_t;wire n4065;wire n4065_t;wire n4066;wire n4066_t;wire n4067;wire n4067_t;wire n4068;wire n4068_t;wire n4069;wire n4069_t;wire n4070;wire n4070_t;wire n4071;wire n4071_t;wire n4072;wire n4072_t;wire n4073;wire n4073_t;wire n4074;wire n4074_t;wire n4075;wire n4075_t;wire n4076;wire n4076_t;wire n4077;wire n4077_t;wire n4078;wire n4078_t;wire n4079;wire n4079_t;wire n4080;wire n4080_t;wire n4081;wire n4081_t;wire n4082;wire n4082_t;wire n4083;wire n4083_t;wire n4084;wire n4084_t;wire n4085;wire n4085_t;wire n4086;wire n4086_t;wire n4087;wire n4087_t;wire n4088;wire n4088_t;wire n4089;wire n4089_t;wire n4090;wire n4090_t;wire n4091;wire n4091_t;wire n4092;wire n4092_t;wire n4093;wire n4093_t;wire n4094;wire n4094_t;wire n4095;wire n4095_t;wire n4096;wire n4096_t;wire n4097;wire n4097_t;wire n4098;wire n4098_t;wire n4099;wire n4099_t;wire n4100;wire n4100_t;wire n4101;wire n4101_t;wire n4102;wire n4102_t;wire n4103;wire n4103_t;wire n4104;wire n4104_t;wire n4105;wire n4105_t;wire n4106;wire n4106_t;wire n4107;wire n4107_t;wire n4108;wire n4108_t;wire n4109;wire n4109_t;wire n4110;wire n4110_t;wire n4111;wire n4111_t;wire n4112;wire n4112_t;wire n4113;wire n4113_t;wire n4114;wire n4114_t;wire n4115;wire n4115_t;wire n4116;wire n4116_t;wire n4117;wire n4117_t;wire n4118;wire n4118_t;wire n4119;wire n4119_t;wire n4120;wire n4120_t;wire n4121;wire n4121_t;wire n4122;wire n4122_t;wire n4123;wire n4123_t;wire n4124;wire n4124_t;wire n4125;wire n4125_t;wire n4126;wire n4126_t;wire n4127;wire n4127_t;wire n4128;wire n4128_t;wire n4129;wire n4129_t;wire n4130;wire n4130_t;wire n4131;wire n4131_t;wire n4132;wire n4132_t;wire n4133;wire n4133_t;wire n4134;wire n4134_t;wire n4135;wire n4135_t;wire n4136;wire n4136_t;wire n4137;wire n4137_t;wire n4138;wire n4138_t;wire n4139;wire n4139_t;wire n4140;wire n4140_t;wire n4141;wire n4141_t;wire n4142;wire n4142_t;wire n4143;wire n4143_t;wire n4144;wire n4144_t;wire n4145;wire n4145_t;wire n4146;wire n4146_t;wire n4147;wire n4147_t;wire n4148;wire n4148_t;wire n4149;wire n4149_t;wire n4150;wire n4150_t;wire n4151;wire n4151_t;wire n4152;wire n4152_t;wire n4153;wire n4153_t;wire n4154;wire n4154_t;wire n4155;wire n4155_t;wire n4156;wire n4156_t;wire n4157;wire n4157_t;wire n4158;wire n4158_t;wire n4159;wire n4159_t;wire n4160;wire n4160_t;wire n4161;wire n4161_t;wire n4162;wire n4162_t;wire n4163;wire n4163_t;wire n4164;wire n4164_t;wire n4165;wire n4165_t;wire n4166;wire n4166_t;wire n4167;wire n4167_t;wire n4168;wire n4168_t;wire n4169;wire n4169_t;wire n4170;wire n4170_t;wire n4171;wire n4171_t;wire n4172;wire n4172_t;wire n4173;wire n4173_t;wire n4174;wire n4174_t;wire n4175;wire n4175_t;wire n4176;wire n4176_t;wire n4177;wire n4177_t;wire n4178;wire n4178_t;wire n4179;wire n4179_t;wire n4180;wire n4180_t;wire n4181;wire n4181_t;wire n4182;wire n4182_t;wire n4183;wire n4183_t;wire n4184;wire n4184_t;wire n4185;wire n4185_t;wire n4186;wire n4186_t;wire n4187;wire n4187_t;wire n4188;wire n4188_t;wire n4189;wire n4189_t;wire n4190;wire n4190_t;wire n4191;wire n4191_t;wire n4192;wire n4192_t;wire n4193;wire n4193_t;wire n4194;wire n4194_t;wire n4195;wire n4195_t;wire n4196;wire n4196_t;wire n4197;wire n4197_t;wire n4198;wire n4198_t;wire n4199;wire n4199_t;wire n4200;wire n4200_t;wire n4201;wire n4201_t;wire n4202;wire n4202_t;wire n4203;wire n4203_t;wire n4204;wire n4204_t;wire n4205;wire n4205_t;wire n4206;wire n4206_t;wire n4207;wire n4207_t;wire n4208;wire n4208_t;wire n4209;wire n4209_t;wire n4210;wire n4210_t;wire n4211;wire n4211_t;wire n4212;wire n4212_t;wire n4213;wire n4213_t;wire n4214;wire n4214_t;wire n4215;wire n4215_t;wire n4216;wire n4216_t;wire n4217;wire n4217_t;wire n4218;wire n4218_t;wire n4219;wire n4219_t;wire n4220;wire n4220_t;wire n4221;wire n4221_t;wire n4222;wire n4222_t;wire n4223;wire n4223_t;wire n4224;wire n4224_t;wire n4225;wire n4225_t;wire n4226;wire n4226_t;wire n4227;wire n4227_t;wire n4228;wire n4228_t;wire n4229;wire n4229_t;wire n4230;wire n4230_t;wire n4231;wire n4231_t;wire n4232;wire n4232_t;wire n4233;wire n4233_t;wire n4234;wire n4234_t;wire n4235;wire n4235_t;wire n4236;wire n4236_t;wire n4237;wire n4237_t;wire n4238;wire n4238_t;wire n4239;wire n4239_t;wire n4240;wire n4240_t;wire n4241;wire n4241_t;wire n4242;wire n4242_t;wire n4243;wire n4243_t;wire n4244;wire n4244_t;wire n4245;wire n4245_t;wire n4246;wire n4246_t;wire n4247;wire n4247_t;wire n4248;wire n4248_t;wire n4249;wire n4249_t;wire n4250;wire n4250_t;wire n4251;wire n4251_t;wire n4252;wire n4252_t;wire n4253;wire n4253_t;wire n4254;wire n4254_t;wire n4255;wire n4255_t;wire n4256;wire n4256_t;wire n4257;wire n4257_t;wire n4258;wire n4258_t;wire n4259;wire n4259_t;wire n4260;wire n4260_t;wire n4261;wire n4261_t;wire n4262;wire n4262_t;wire n4263;wire n4263_t;wire n4264;wire n4264_t;wire n4265;wire n4265_t;wire n4266;wire n4266_t;wire n4267;wire n4267_t;wire n4268;wire n4268_t;wire n4269;wire n4269_t;wire n4270;wire n4270_t;wire n4271;wire n4271_t;wire n4272;wire n4272_t;wire n4273;wire n4273_t;wire n4274;wire n4274_t;wire n4275;wire n4275_t;wire n4276;wire n4276_t;wire n4277;wire n4277_t;wire n4278;wire n4278_t;wire n4279;wire n4279_t;wire n4280;wire n4280_t;wire n4281;wire n4281_t;wire n4282;wire n4282_t;wire n4283;wire n4283_t;wire n4284;wire n4284_t;wire n4285;wire n4285_t;wire n4286;wire n4286_t;wire n4287;wire n4287_t;wire n4288;wire n4288_t;wire n4289;wire n4289_t;wire n4290;wire n4290_t;wire n4291;wire n4291_t;wire n4292;wire n4292_t;wire n4293;wire n4293_t;wire n4294;wire n4294_t;wire n4295;wire n4295_t;wire n4296;wire n4296_t;wire n4297;wire n4297_t;wire n4298;wire n4298_t;wire n4299;wire n4299_t;wire n4300;wire n4300_t;wire n4301;wire n4301_t;wire n4302;wire n4302_t;wire n4303;wire n4303_t;wire n4304;wire n4304_t;wire n4305;wire n4305_t;wire n4306;wire n4306_t;wire n4307;wire n4307_t;wire n4308;wire n4308_t;wire n4309;wire n4309_t;wire n4310;wire n4310_t;wire n4311;wire n4311_t;wire n4312;wire n4312_t;wire n4313;wire n4313_t;wire n4314;wire n4314_t;wire n4315;wire n4315_t;wire n4316;wire n4316_t;wire n4317;wire n4317_t;wire n4318;wire n4318_t;wire n4319;wire n4319_t;wire n4320;wire n4320_t;wire n4321;wire n4321_t;wire n4322;wire n4322_t;wire n4323;wire n4323_t;wire n4324;wire n4324_t;wire n4325;wire n4325_t;wire n4326;wire n4326_t;wire n4327;wire n4327_t;wire n4328;wire n4328_t;wire n4329;wire n4329_t;wire n4330;wire n4330_t;wire n4331;wire n4331_t;wire n4332;wire n4332_t;wire n4333;wire n4333_t;wire n4334;wire n4334_t;wire n4335;wire n4335_t;wire n4336;wire n4336_t;wire n4337;wire n4337_t;wire n4338;wire n4338_t;wire n4339;wire n4339_t;wire n4340;wire n4340_t;wire n4341;wire n4341_t;wire n4342;wire n4342_t;wire n4343;wire n4343_t;wire n4344;wire n4344_t;wire n4345;wire n4345_t;wire n4346;wire n4346_t;wire n4347;wire n4347_t;wire n4348;wire n4348_t;wire n4349;wire n4349_t;wire n4350;wire n4350_t;wire n4351;wire n4351_t;wire n4352;wire n4352_t;wire n4353;wire n4353_t;wire n4354;wire n4354_t;wire n4355;wire n4355_t;wire n4356;wire n4356_t;wire n4357;wire n4357_t;wire n4358;wire n4358_t;wire n4359;wire n4359_t;wire n4360;wire n4360_t;wire n4361;wire n4361_t;wire n4362;wire n4362_t;wire n4363;wire n4363_t;wire n4364;wire n4364_t;wire n4365;wire n4365_t;wire n4366;wire n4366_t;wire n4367;wire n4367_t;wire n4368;wire n4368_t;wire n4369;wire n4369_t;wire n4370;wire n4370_t;wire n4371;wire n4371_t;wire n4372;wire n4372_t;wire n4373;wire n4373_t;wire n4374;wire n4374_t;wire n4375;wire n4375_t;wire n4376;wire n4376_t;wire n4377;wire n4377_t;wire n4378;wire n4378_t;wire n4379;wire n4379_t;wire n4380;wire n4380_t;wire n4381;wire n4381_t;wire n4382;wire n4382_t;wire n4383;wire n4383_t;wire n4384;wire n4384_t;wire n4385;wire n4385_t;wire n4386;wire n4386_t;wire n4387;wire n4387_t;wire n4388;wire n4388_t;wire n4389;wire n4389_t;wire n4390;wire n4390_t;wire n4391;wire n4391_t;wire n4392;wire n4392_t;wire n4393;wire n4393_t;wire n4394;wire n4394_t;wire n4395;wire n4395_t;wire n4396;wire n4396_t;wire n4397;wire n4397_t;wire n4398;wire n4398_t;wire n4399;wire n4399_t;wire n4400;wire n4400_t;wire n4401;wire n4401_t;wire n4402;wire n4402_t;wire n4403;wire n4403_t;wire n4404;wire n4404_t;wire n4405;wire n4405_t;wire n4406;wire n4406_t;wire n4407;wire n4407_t;wire n4408;wire n4408_t;wire n4409;wire n4409_t;wire n4410;wire n4410_t;wire n4411;wire n4411_t;wire n4412;wire n4412_t;wire n4413;wire n4413_t;wire n4414;wire n4414_t;wire n4415;wire n4415_t;wire n4416;wire n4416_t;wire n4417;wire n4417_t;wire n4418;wire n4418_t;wire n4419;wire n4419_t;wire n4420;wire n4420_t;wire n4421;wire n4421_t;wire n4422;wire n4422_t;wire n4423;wire n4423_t;wire n4424;wire n4424_t;wire n4425;wire n4425_t;wire n4426;wire n4426_t;wire n4427;wire n4427_t;wire n4428;wire n4428_t;wire n4429;wire n4429_t;wire n4430;wire n4430_t;wire n4431;wire n4431_t;wire n4432;wire n4432_t;wire n4433;wire n4433_t;wire n4434;wire n4434_t;wire n4435;wire n4435_t;wire n4436;wire n4436_t;wire n4437;wire n4437_t;wire n4438;wire n4438_t;wire n4439;wire n4439_t;wire n4440;wire n4440_t;wire n4441;wire n4441_t;wire n4442;wire n4442_t;wire n4443;wire n4443_t;wire n4444;wire n4444_t;wire n4445;wire n4445_t;wire n4446;wire n4446_t;wire n4447;wire n4447_t;wire n4448;wire n4448_t;wire n4449;wire n4449_t;wire n4450;wire n4450_t;wire n4451;wire n4451_t;wire n4452;wire n4452_t;wire n4453;wire n4453_t;wire n4454;wire n4454_t;wire n4455;wire n4455_t;wire n4456;wire n4456_t;wire n4457;wire n4457_t;wire n4458;wire n4458_t;wire n4459;wire n4459_t;wire n4460;wire n4460_t;wire n4461;wire n4461_t;wire n4462;wire n4462_t;wire n4463;wire n4463_t;wire n4464;wire n4464_t;wire n4465;wire n4465_t;wire n4466;wire n4466_t;wire n4467;wire n4467_t;wire n4468;wire n4468_t;wire n4469;wire n4469_t;wire n4470;wire n4470_t;wire n4471;wire n4471_t;wire n4472;wire n4472_t;wire n4473;wire n4473_t;wire n4474;wire n4474_t;wire n4475;wire n4475_t;wire n4476;wire n4476_t;wire n4477;wire n4477_t;wire n4478;wire n4478_t;wire n4479;wire n4479_t;wire n4480;wire n4480_t;wire n4481;wire n4481_t;wire n4482;wire n4482_t;wire n4483;wire n4483_t;wire n4484;wire n4484_t;wire n4485;wire n4485_t;wire n4486;wire n4486_t;wire n4487;wire n4487_t;wire n4488;wire n4488_t;wire n4489;wire n4489_t;wire n4490;wire n4490_t;wire n4491;wire n4491_t;wire n4492;wire n4492_t;wire n4493;wire n4493_t;wire n4494;wire n4494_t;wire n4495;wire n4495_t;wire n4496;wire n4496_t;wire n4497;wire n4497_t;wire n4498;wire n4498_t;wire n4499;wire n4499_t;wire n4500;wire n4500_t;wire n4501;wire n4501_t;wire n4502;wire n4502_t;wire n4503;wire n4503_t;wire n4504;wire n4504_t;wire n4505;wire n4505_t;wire n4506;wire n4506_t;wire n4507;wire n4507_t;wire n4508;wire n4508_t;wire n4509;wire n4509_t;wire n4510;wire n4510_t;wire n4511;wire n4511_t;wire n4512;wire n4512_t;wire n4513;wire n4513_t;wire n4514;wire n4514_t;wire n4515;wire n4515_t;wire n4516;wire n4516_t;wire n4517;wire n4517_t;wire n4518;wire n4518_t;wire n4519;wire n4519_t;wire n4520;wire n4520_t;wire n4521;wire n4521_t;wire n4522;wire n4522_t;wire n4523;wire n4523_t;wire n4524;wire n4524_t;wire n4525;wire n4525_t;wire n4526;wire n4526_t;wire n4527;wire n4527_t;wire n4528;wire n4528_t;wire n4529;wire n4529_t;wire n4530;wire n4530_t;wire n4531;wire n4531_t;wire n4532;wire n4532_t;wire n4533;wire n4533_t;wire n4534;wire n4534_t;wire n4535;wire n4535_t;wire n4536;wire n4536_t;wire n4537;wire n4537_t;wire n4538;wire n4538_t;wire n4539;wire n4539_t;wire n4540;wire n4540_t;wire n4541;wire n4541_t;wire n4542;wire n4542_t;wire n4543;wire n4543_t;wire n4544;wire n4544_t;wire n4545;wire n4545_t;wire n4546;wire n4546_t;wire n4547;wire n4547_t;wire n4548;wire n4548_t;wire n4549;wire n4549_t;wire n4550;wire n4550_t;wire n4551;wire n4551_t;wire n4552;wire n4552_t;wire n4553;wire n4553_t;wire n4554;wire n4554_t;wire n4555;wire n4555_t;wire n4556;wire n4556_t;wire n4557;wire n4557_t;wire n4558;wire n4558_t;wire n4559;wire n4559_t;wire n4560;wire n4560_t;wire n4561;wire n4561_t;wire n4562;wire n4562_t;wire n4563;wire n4563_t;wire n4564;wire n4564_t;wire n4565;wire n4565_t;wire n4566;wire n4566_t;wire n4567;wire n4567_t;wire n4568;wire n4568_t;wire n4569;wire n4569_t;wire n4570;wire n4570_t;wire n4571;wire n4571_t;wire n4572;wire n4572_t;wire n4573;wire n4573_t;wire n4574;wire n4574_t;wire n4575;wire n4575_t;wire n4576;wire n4576_t;wire n4577;wire n4577_t;wire n4578;wire n4578_t;wire n4579;wire n4579_t;wire n4580;wire n4580_t;wire n4581;wire n4581_t;wire n4582;wire n4582_t;wire n4583;wire n4583_t;wire n4584;wire n4584_t;wire n4585;wire n4585_t;wire n4586;wire n4586_t;wire n4587;wire n4587_t;wire n4588;wire n4588_t;wire n4589;wire n4589_t;wire n4590;wire n4590_t;wire n4591;wire n4591_t;wire n4592;wire n4592_t;wire n4593;wire n4593_t;wire n4594;wire n4594_t;wire n4595;wire n4595_t;wire n4596;wire n4596_t;wire n4597;wire n4597_t;wire n4598;wire n4598_t;wire n4599;wire n4599_t;wire n4600;wire n4600_t;wire n4601;wire n4601_t;wire n4602;wire n4602_t;wire n4603;wire n4603_t;wire n4604;wire n4604_t;wire n4605;wire n4605_t;wire n4606;wire n4606_t;wire n4607;wire n4607_t;wire n4608;wire n4608_t;wire n4609;wire n4609_t;wire n4610;wire n4610_t;wire n4611;wire n4611_t;wire n4612;wire n4612_t;wire n4613;wire n4613_t;wire n4614;wire n4614_t;wire n4615;wire n4615_t;wire n4616;wire n4616_t;wire n4617;wire n4617_t;wire n4618;wire n4618_t;wire n4619;wire n4619_t;wire n4620;wire n4620_t;wire n4621;wire n4621_t;wire n4622;wire n4622_t;wire n4623;wire n4623_t;wire n4624;wire n4624_t;wire n4625;wire n4625_t;wire n4626;wire n4626_t;wire n4627;wire n4627_t;wire n4628;wire n4628_t;wire n4629;wire n4629_t;wire n4630;wire n4630_t;wire n4631;wire n4631_t;wire n4632;wire n4632_t;wire n4633;wire n4633_t;wire n4634;wire n4634_t;wire n4635;wire n4635_t;wire n4636;wire n4636_t;wire n4637;wire n4637_t;wire n4638;wire n4638_t;wire n4639;wire n4639_t;wire n4640;wire n4640_t;wire n4641;wire n4641_t;wire n4642;wire n4642_t;wire n4643;wire n4643_t;wire n4644;wire n4644_t;wire n4645;wire n4645_t;wire n4646;wire n4646_t;wire n4647;wire n4647_t;wire n4648;wire n4648_t;wire n4649;wire n4649_t;wire n4650;wire n4650_t;wire n4651;wire n4651_t;wire n4652;wire n4652_t;wire n4653;wire n4653_t;wire n4654;wire n4654_t;wire n4655;wire n4655_t;wire n4656;wire n4656_t;wire n4657;wire n4657_t;wire n4658;wire n4658_t;wire n4659;wire n4659_t;wire n4660;wire n4660_t;wire n4661;wire n4661_t;wire n4662;wire n4662_t;wire n4663;wire n4663_t;wire n4664;wire n4664_t;wire n4665;wire n4665_t;wire n4666;wire n4666_t;wire n4667;wire n4667_t;wire n4668;wire n4668_t;wire n4669;wire n4669_t;wire n4670;wire n4670_t;wire n4671;wire n4671_t;wire n4672;wire n4672_t;wire n4673;wire n4673_t;wire n4674;wire n4674_t;wire n4675;wire n4675_t;wire n4676;wire n4676_t;wire n4677;wire n4677_t;wire n4678;wire n4678_t;wire n4679;wire n4679_t;wire n4680;wire n4680_t;wire n4681;wire n4681_t;wire n4682;wire n4682_t;wire n4683;wire n4683_t;wire n4684;wire n4684_t;wire n4685;wire n4685_t;wire n4686;wire n4686_t;wire n4687;wire n4687_t;wire n4688;wire n4688_t;wire n4689;wire n4689_t;wire n4690;wire n4690_t;wire n4691;wire n4691_t;wire n4692;wire n4692_t;wire n4693;wire n4693_t;wire n4694;wire n4694_t;wire n4695;wire n4695_t;wire n4696;wire n4696_t;wire n4697;wire n4697_t;wire n4698;wire n4698_t;wire n4699;wire n4699_t;wire n4700;wire n4700_t;wire n4701;wire n4701_t;wire n4702;wire n4702_t;wire n4703;wire n4703_t;wire n4704;wire n4704_t;wire n4705;wire n4705_t;wire n4706;wire n4706_t;wire n4707;wire n4707_t;wire n4708;wire n4708_t;wire n4709;wire n4709_t;wire n4710;wire n4710_t;wire n4711;wire n4711_t;wire n4712;wire n4712_t;wire n4713;wire n4713_t;wire n4714;wire n4714_t;wire n4715;wire n4715_t;wire n4716;wire n4716_t;wire n4717;wire n4717_t;wire n4718;wire n4718_t;wire n4719;wire n4719_t;wire n4720;wire n4720_t;wire n4721;wire n4721_t;wire n4722;wire n4722_t;wire n4723;wire n4723_t;wire n4724;wire n4724_t;wire n4725;wire n4725_t;wire n4726;wire n4726_t;wire n4727;wire n4727_t;wire n4728;wire n4728_t;wire n4729;wire n4729_t;wire n4730;wire n4730_t;wire n4731;wire n4731_t;wire n4732;wire n4732_t;wire n4733;wire n4733_t;wire n4734;wire n4734_t;wire n4735;wire n4735_t;wire n4736;wire n4736_t;wire n4737;wire n4737_t;wire n4738;wire n4738_t;wire n4739;wire n4739_t;wire n4740;wire n4740_t;wire n4741;wire n4741_t;wire n4742;wire n4742_t;wire n4743;wire n4743_t;wire n4744;wire n4744_t;wire n4745;wire n4745_t;wire n4746;wire n4746_t;wire n4747;wire n4747_t;wire n4748;wire n4748_t;wire n4749;wire n4749_t;wire n4750;wire n4750_t;wire n4751;wire n4751_t;wire n4752;wire n4752_t;wire n4753;wire n4753_t;wire n4754;wire n4754_t;wire n4755;wire n4755_t;wire n4756;wire n4756_t;wire n4757;wire n4757_t;wire n4758;wire n4758_t;wire n4759;wire n4759_t;wire n4760;wire n4760_t;wire n4761;wire n4761_t;wire n4762;wire n4762_t;wire n4763;wire n4763_t;wire n4764;wire n4764_t;wire n4765;wire n4765_t;wire n4766;wire n4766_t;wire n4767;wire n4767_t;wire n4768;wire n4768_t;wire n4769;wire n4769_t;wire n4770;wire n4770_t;wire n4771;wire n4771_t;wire n4772;wire n4772_t;wire n4773;wire n4773_t;wire n4774;wire n4774_t;wire n4775;wire n4775_t;wire n4776;wire n4776_t;wire n4777;wire n4777_t;wire n4778;wire n4778_t;wire n4779;wire n4779_t;wire n4780;wire n4780_t;wire n4781;wire n4781_t;wire n4782;wire n4782_t;wire n4783;wire n4783_t;wire n4784;wire n4784_t;wire n4785;wire n4785_t;wire n4786;wire n4786_t;wire n4787;wire n4787_t;wire n4788;wire n4788_t;wire n4789;wire n4789_t;wire n4790;wire n4790_t;wire n4791;wire n4791_t;wire n4792;wire n4792_t;wire n4793;wire n4793_t;wire n4794;wire n4794_t;wire n4795;wire n4795_t;wire n4796;wire n4796_t;wire n4797;wire n4797_t;wire n4798;wire n4798_t;wire n4799;wire n4799_t;wire n4800;wire n4800_t;wire n4801;wire n4801_t;wire n4802;wire n4802_t;wire n4803;wire n4803_t;wire n4804;wire n4804_t;wire n4805;wire n4805_t;wire n4806;wire n4806_t;wire n4807;wire n4807_t;wire n4808;wire n4808_t;wire n4809;wire n4809_t;wire n4810;wire n4810_t;wire n4811;wire n4811_t;wire n4812;wire n4812_t;wire n4813;wire n4813_t;wire n4814;wire n4814_t;wire n4815;wire n4815_t;wire n4816;wire n4816_t;wire n4817;wire n4817_t;wire n4818;wire n4818_t;wire n4819;wire n4819_t;wire n4820;wire n4820_t;wire n4821;wire n4821_t;wire n4822;wire n4822_t;wire n4823;wire n4823_t;wire n4824;wire n4824_t;wire n4825;wire n4825_t;wire n4826;wire n4826_t;wire n4827;wire n4827_t;wire n4828;wire n4828_t;wire n4829;wire n4829_t;wire n4830;wire n4830_t;wire n4831;wire n4831_t;wire n4832;wire n4832_t;wire n4833;wire n4833_t;wire n4834;wire n4834_t;wire n4835;wire n4835_t;wire n4836;wire n4836_t;wire n4837;wire n4837_t;wire n4838;wire n4838_t;wire n4839;wire n4839_t;wire n4840;wire n4840_t;wire n4841;wire n4841_t;wire n4842;wire n4842_t;wire n4843;wire n4843_t;wire n4844;wire n4844_t;wire n4845;wire n4845_t;wire n4846;wire n4846_t;wire n4847;wire n4847_t;wire n4848;wire n4848_t;wire n4849;wire n4849_t;wire n4850;wire n4850_t;wire n4851;wire n4851_t;wire n4852;wire n4852_t;wire n4853;wire n4853_t;wire n4854;wire n4854_t;wire n4855;wire n4855_t;wire n4856;wire n4856_t;wire n4857;wire n4857_t;wire n4858;wire n4858_t;wire n4859;wire n4859_t;wire n4860;wire n4860_t;wire n4861;wire n4861_t;wire n4862;wire n4862_t;wire n4863;wire n4863_t;wire n4864;wire n4864_t;wire n4865;wire n4865_t;wire n4866;wire n4866_t;wire n4867;wire n4867_t;wire n4868;wire n4868_t;wire n4869;wire n4869_t;wire n4870;wire n4870_t;wire n4871;wire n4871_t;wire n4872;wire n4872_t;wire n4873;wire n4873_t;wire n4874;wire n4874_t;wire n4875;wire n4875_t;wire n4876;wire n4876_t;wire n4877;wire n4877_t;wire n4878;wire n4878_t;wire n4879;wire n4879_t;wire n4880;wire n4880_t;wire n4881;wire n4881_t;wire n4882;wire n4882_t;wire n4883;wire n4883_t;wire n4884;wire n4884_t;wire n4885;wire n4885_t;wire n4886;wire n4886_t;wire n4887;wire n4887_t;wire n4888;wire n4888_t;wire n4889;wire n4889_t;wire n4890;wire n4890_t;wire n4891;wire n4891_t;wire n4892;wire n4892_t;wire n4893;wire n4893_t;wire n4894;wire n4894_t;wire n4895;wire n4895_t;wire n4896;wire n4896_t;wire n4897;wire n4897_t;wire n4898;wire n4898_t;wire n4899;wire n4899_t;wire n4900;wire n4900_t;wire n4901;wire n4901_t;wire n4902;wire n4902_t;wire n4903;wire n4903_t;wire n4904;wire n4904_t;wire n4905;wire n4905_t;wire n4906;wire n4906_t;wire n4907;wire n4907_t;wire n4908;wire n4908_t;wire n4909;wire n4909_t;wire n4910;wire n4910_t;wire n4911;wire n4911_t;wire n4912;wire n4912_t;wire n4913;wire n4913_t;wire n4914;wire n4914_t;wire n4915;wire n4915_t;wire n4916;wire n4916_t;wire n4917;wire n4917_t;wire n4918;wire n4918_t;wire n4919;wire n4919_t;wire n4920;wire n4920_t;wire n4921;wire n4921_t;wire n4922;wire n4922_t;wire n4923;wire n4923_t;wire n4924;wire n4924_t;wire n4925;wire n4925_t;wire n4926;wire n4926_t;wire n4927;wire n4927_t;wire n4928;wire n4928_t;wire n4929;wire n4929_t;wire n4930;wire n4930_t;wire n4931;wire n4931_t;wire n4932;wire n4932_t;wire n4933;wire n4933_t;wire n4934;wire n4934_t;wire n4935;wire n4935_t;wire n4936;wire n4936_t;wire n4937;wire n4937_t;wire n4938;wire n4938_t;wire n4939;wire n4939_t;wire n4940;wire n4940_t;wire n4941;wire n4941_t;wire n4942;wire n4942_t;wire n4943;wire n4943_t;wire n4944;wire n4944_t;wire n4945;wire n4945_t;wire n4946;wire n4946_t;wire n4947;wire n4947_t;wire n4948;wire n4948_t;wire n4949;wire n4949_t;wire n4950;wire n4950_t;wire n4951;wire n4951_t;wire n4952;wire n4952_t;wire n4953;wire n4953_t;wire n4954;wire n4954_t;wire n4955;wire n4955_t;wire n4956;wire n4956_t;wire n4957;wire n4957_t;wire n4958;wire n4958_t;wire n4959;wire n4959_t;wire n4960;wire n4960_t;wire n4961;wire n4961_t;wire n4962;wire n4962_t;wire n4963;wire n4963_t;wire n4964;wire n4964_t;wire n4965;wire n4965_t;wire n4966;wire n4966_t;wire n4967;wire n4967_t;wire n4968;wire n4968_t;wire n4969;wire n4969_t;wire n4970;wire n4970_t;wire n4971;wire n4971_t;wire n4972;wire n4972_t;wire n4973;wire n4973_t;wire n4974;wire n4974_t;wire n4975;wire n4975_t;wire n4976;wire n4976_t;wire n4977;wire n4977_t;wire n4978;wire n4978_t;wire n4979;wire n4979_t;wire n4980;wire n4980_t;wire n4981;wire n4981_t;wire n4982;wire n4982_t;wire n4983;wire n4983_t;wire n4984;wire n4984_t;wire n4985;wire n4985_t;wire n4986;wire n4986_t;wire n4987;wire n4987_t;wire n4988;wire n4988_t;wire n4989;wire n4989_t;wire n4990;wire n4990_t;wire n4991;wire n4991_t;wire n4992;wire n4992_t;wire n4993;wire n4993_t;wire n4994;wire n4994_t;wire n4995;wire n4995_t;wire n4996;wire n4996_t;wire n4997;wire n4997_t;wire n4998;wire n4998_t;wire n4999;wire n4999_t;wire n5000;wire n5000_t;wire n5001;wire n5001_t;wire n5002;wire n5002_t;wire n5003;wire n5003_t;wire n5004;wire n5004_t;wire n5005;wire n5005_t;wire n5006;wire n5006_t;wire n5007;wire n5007_t;wire n5008;wire n5008_t;wire n5009;wire n5009_t;wire n5010;wire n5010_t;wire n5011;wire n5011_t;wire n5012;wire n5012_t;wire n5013;wire n5013_t;wire n5014;wire n5014_t;wire n5015;wire n5015_t;wire n5016;wire n5016_t;wire n5017;wire n5017_t;wire n5018;wire n5018_t;wire n5019;wire n5019_t;wire n5020;wire n5020_t;wire n5021;wire n5021_t;wire n5022;wire n5022_t;wire n5023;wire n5023_t;wire n5024;wire n5024_t;wire n5025;wire n5025_t;wire n5026;wire n5026_t;wire n5027;wire n5027_t;wire n5028;wire n5028_t;wire n5029;wire n5029_t;wire n5030;wire n5030_t;wire n5031;wire n5031_t;wire n5032;wire n5032_t;wire n5033;wire n5033_t;wire n5034;wire n5034_t;wire n5035;wire n5035_t;wire n5036;wire n5036_t;wire n5037;wire n5037_t;wire n5038;wire n5038_t;wire n5039;wire n5039_t;wire n5040;wire n5040_t;wire n5041;wire n5041_t;wire n5042;wire n5042_t;wire n5043;wire n5043_t;wire n5044;wire n5044_t;wire n5045;wire n5045_t;wire n5046;wire n5046_t;wire n5047;wire n5047_t;wire n5048;wire n5048_t;wire n5049;wire n5049_t;wire n5050;wire n5050_t;wire n5051;wire n5051_t;wire n5052;wire n5052_t;wire n5053;wire n5053_t;wire n5054;wire n5054_t;wire n5055;wire n5055_t;wire n5056;wire n5056_t;wire n5057;wire n5057_t;wire n5058;wire n5058_t;wire n5059;wire n5059_t;wire n5060;wire n5060_t;wire n5061;wire n5061_t;wire n5062;wire n5062_t;wire n5063;wire n5063_t;wire n5064;wire n5064_t;wire n5065;wire n5065_t;wire n5066;wire n5066_t;wire n5067;wire n5067_t;wire n5068;wire n5068_t;wire n5069;wire n5069_t;wire n5070;wire n5070_t;wire n5071;wire n5071_t;wire n5072;wire n5072_t;wire n5073;wire n5073_t;wire n5074;wire n5074_t;wire n5075;wire n5075_t;wire n5076;wire n5076_t;wire n5077;wire n5077_t;wire n5078;wire n5078_t;wire n5079;wire n5079_t;wire n5080;wire n5080_t;wire n5081;wire n5081_t;wire n5082;wire n5082_t;wire n5083;wire n5083_t;wire n5084;wire n5084_t;wire n5085;wire n5085_t;wire n5086;wire n5086_t;wire n5087;wire n5087_t;wire n5088;wire n5088_t;wire n5089;wire n5089_t;wire n5090;wire n5090_t;wire n5091;wire n5091_t;wire n5092;wire n5092_t;wire n5093;wire n5093_t;wire n5094;wire n5094_t;wire n5095;wire n5095_t;wire n5096;wire n5096_t;wire n5097;wire n5097_t;wire n5098;wire n5098_t;wire n5099;wire n5099_t;wire n5100;wire n5100_t;wire n5101;wire n5101_t;wire n5102;wire n5102_t;wire n5103;wire n5103_t;wire n5104;wire n5104_t;wire n5105;wire n5105_t;wire n5106;wire n5106_t;wire n5107;wire n5107_t;wire n5108;wire n5108_t;wire n5109;wire n5109_t;wire n5110;wire n5110_t;wire n5111;wire n5111_t;wire n5112;wire n5112_t;wire n5113;wire n5113_t;wire n5114;wire n5114_t;wire n5115;wire n5115_t;wire n5116;wire n5116_t;wire n5117;wire n5117_t;wire n5118;wire n5118_t;wire n5119;wire n5119_t;wire n5120;wire n5120_t;wire n5121;wire n5121_t;wire n5122;wire n5122_t;wire n5123;wire n5123_t;wire n5124;wire n5124_t;wire n5125;wire n5125_t;wire n5126;wire n5126_t;wire n5127;wire n5127_t;wire n5128;wire n5128_t;wire n5129;wire n5129_t;wire n5130;wire n5130_t;wire n5131;wire n5131_t;wire n5132;wire n5132_t;wire n5133;wire n5133_t;wire n5134;wire n5134_t;wire n5135;wire n5135_t;wire n5136;wire n5136_t;wire n5137;wire n5137_t;wire n5138;wire n5138_t;wire n5139;wire n5139_t;wire n5140;wire n5140_t;wire n5141;wire n5141_t;wire n5142;wire n5142_t;wire n5143;wire n5143_t;wire n5144;wire n5144_t;wire n5145;wire n5145_t;wire n5146;wire n5146_t;wire n5147;wire n5147_t;wire n5148;wire n5148_t;wire n5149;wire n5149_t;wire n5150;wire n5150_t;wire n5151;wire n5151_t;wire n5152;wire n5152_t;wire n5153;wire n5153_t;wire n5154;wire n5154_t;wire n5155;wire n5155_t;wire n5156;wire n5156_t;wire n5157;wire n5157_t;wire n5158;wire n5158_t;wire n5159;wire n5159_t;wire n5160;wire n5160_t;wire n5161;wire n5161_t;wire n5162;wire n5162_t;wire n5163;wire n5163_t;wire n5164;wire n5164_t;wire n5165;wire n5165_t;wire n5166;wire n5166_t;wire n5167;wire n5167_t;wire n5168;wire n5168_t;wire n5169;wire n5169_t;wire n5170;wire n5170_t;wire n5171;wire n5171_t;wire n5172;wire n5172_t;wire n5173;wire n5173_t;wire n5174;wire n5174_t;wire n5175;wire n5175_t;wire n5176;wire n5176_t;wire n5177;wire n5177_t;wire n5178;wire n5178_t;wire n5179;wire n5179_t;wire n5180;wire n5180_t;wire n5181;wire n5181_t;wire n5182;wire n5182_t;wire n5183;wire n5183_t;wire n5184;wire n5184_t;wire n5185;wire n5185_t;wire n5186;wire n5186_t;wire n5187;wire n5187_t;wire n5188;wire n5188_t;wire n5189;wire n5189_t;wire n5190;wire n5190_t;wire n5191;wire n5191_t;wire n5192;wire n5192_t;wire n5193;wire n5193_t;wire n5194;wire n5194_t;wire n5195;wire n5195_t;wire n5196;wire n5196_t;wire n5197;wire n5197_t;wire n5198;wire n5198_t;wire n5199;wire n5199_t;wire n5200;wire n5200_t;wire n5201;wire n5201_t;wire n5202;wire n5202_t;wire n5203;wire n5203_t;wire n5204;wire n5204_t;wire n5205;wire n5205_t;wire n5206;wire n5206_t;wire n5207;wire n5207_t;wire n5208;wire n5208_t;wire n5209;wire n5209_t;wire n5210;wire n5210_t;wire n5211;wire n5211_t;wire n5212;wire n5212_t;wire n5213;wire n5213_t;wire n5214;wire n5214_t;wire n5215;wire n5215_t;wire n5216;wire n5216_t;wire n5217;wire n5217_t;wire n5218;wire n5218_t;wire n5219;wire n5219_t;wire n5220;wire n5220_t;wire n5221;wire n5221_t;wire n5222;wire n5222_t;wire n5223;wire n5223_t;wire n5224;wire n5224_t;wire n5225;wire n5225_t;wire n5226;wire n5226_t;wire n5227;wire n5227_t;wire n5228;wire n5228_t;wire n5229;wire n5229_t;wire n5230;wire n5230_t;wire n5231;wire n5231_t;wire n5232;wire n5232_t;wire n5233;wire n5233_t;wire n5234;wire n5234_t;wire n5235;wire n5235_t;wire n5236;wire n5236_t;wire n5237;wire n5237_t;wire n5238;wire n5238_t;wire n5239;wire n5239_t;wire n5240;wire n5240_t;wire n5241;wire n5241_t;wire n5242;wire n5242_t;wire n5243;wire n5243_t;wire n5244;wire n5244_t;wire n5245;wire n5245_t;wire n5246;wire n5246_t;wire n5247;wire n5247_t;wire n5248;wire n5248_t;wire n5249;wire n5249_t;wire n5250;wire n5250_t;wire n5251;wire n5251_t;wire n5252;wire n5252_t;wire n5253;wire n5253_t;wire n5254;wire n5254_t;wire n5255;wire n5255_t;wire n5256;wire n5256_t;wire n5257;wire n5257_t;wire n5258;wire n5258_t;wire n5259;wire n5259_t;wire n5260;wire n5260_t;wire n5261;wire n5261_t;wire n5262;wire n5262_t;wire n5263;wire n5263_t;wire n5264;wire n5264_t;wire n5265;wire n5265_t;wire n5266;wire n5266_t;wire n5267;wire n5267_t;wire n5268;wire n5268_t;wire n5269;wire n5269_t;wire n5270;wire n5270_t;wire n5271;wire n5271_t;wire n5272;wire n5272_t;wire n5273;wire n5273_t;wire n5274;wire n5274_t;wire n5275;wire n5275_t;wire n5276;wire n5276_t;wire n5277;wire n5277_t;wire n5278;wire n5278_t;wire n5279;wire n5279_t;wire n5280;wire n5280_t;wire n5281;wire n5281_t;wire n5282;wire n5282_t;wire n5283;wire n5283_t;wire n5284;wire n5284_t;wire n5285;wire n5285_t;wire n5286;wire n5286_t;wire n5287;wire n5287_t;wire n5288;wire n5288_t;wire n5289;wire n5289_t;wire n5290;wire n5290_t;wire n5291;wire n5291_t;wire n5292;wire n5292_t;wire n5293;wire n5293_t;wire n5294;wire n5294_t;wire n5295;wire n5295_t;wire n5296;wire n5296_t;wire n5297;wire n5297_t;wire n5298;wire n5298_t;wire n5299;wire n5299_t;wire n5300;wire n5300_t;wire n5301;wire n5301_t;wire n5302;wire n5302_t;wire n5303;wire n5303_t;wire n5304;wire n5304_t;wire n5305;wire n5305_t;wire n5306;wire n5306_t;wire n5307;wire n5307_t;wire n5308;wire n5308_t;wire n5309;wire n5309_t;wire n5310;wire n5310_t;wire n5311;wire n5311_t;wire n5312;wire n5312_t;wire n5313;wire n5313_t;wire n5314;wire n5314_t;wire n5315;wire n5315_t;wire n5316;wire n5316_t;wire n5317;wire n5317_t;wire n5318;wire n5318_t;wire n5319;wire n5319_t;wire n5320;wire n5320_t;wire n5321;wire n5321_t;wire n5322;wire n5322_t;wire n5323;wire n5323_t;wire n5324;wire n5324_t;wire n5325;wire n5325_t;wire n5326;wire n5326_t;wire n5327;wire n5327_t;wire n5328;wire n5328_t;wire n5329;wire n5329_t;wire n5330;wire n5330_t;wire n5331;wire n5331_t;wire n5332;wire n5332_t;wire n5333;wire n5333_t;wire n5334;wire n5334_t;wire n5335;wire n5335_t;wire n5336;wire n5336_t;wire n5337;wire n5337_t;wire n5338;wire n5338_t;wire n5339;wire n5339_t;wire n5340;wire n5340_t;wire n5341;wire n5341_t;wire n5342;wire n5342_t;wire n5343;wire n5343_t;wire n5344;wire n5344_t;wire n5345;wire n5345_t;wire n5346;wire n5346_t;wire n5347;wire n5347_t;wire n5348;wire n5348_t;wire n5349;wire n5349_t;wire n5350;wire n5350_t;wire n5351;wire n5351_t;wire n5352;wire n5352_t;wire n5353;wire n5353_t;wire n5354;wire n5354_t;wire n5355;wire n5355_t;wire n5356;wire n5356_t;wire n5357;wire n5357_t;wire n5358;wire n5358_t;wire n5359;wire n5359_t;wire n5360;wire n5360_t;wire n5361;wire n5361_t;wire n5362;wire n5362_t;wire n5363;wire n5363_t;wire n5364;wire n5364_t;wire n5365;wire n5365_t;wire n5366;wire n5366_t;wire n5367;wire n5367_t;wire n5368;wire n5368_t;wire n5369;wire n5369_t;wire n5370;wire n5370_t;wire n5371;wire n5371_t;wire n5372;wire n5372_t;wire n5373;wire n5373_t;wire n5374;wire n5374_t;wire n5375;wire n5375_t;wire n5376;wire n5376_t;wire n5377;wire n5377_t;wire n5378;wire n5378_t;wire n5379;wire n5379_t;wire n5380;wire n5380_t;wire n5381;wire n5381_t;wire n5382;wire n5382_t;wire n5383;wire n5383_t;wire n5384;wire n5384_t;wire n5385;wire n5385_t;wire n5386;wire n5386_t;wire n5387;wire n5387_t;wire n5388;wire n5388_t;wire n5389;wire n5389_t;wire n5390;wire n5390_t;wire n5391;wire n5391_t;wire n5392;wire n5392_t;wire n5393;wire n5393_t;wire n5394;wire n5394_t;wire n5395;wire n5395_t;wire n5396;wire n5396_t;wire n5397;wire n5397_t;wire n5398;wire n5398_t;wire n5399;wire n5399_t;wire n5400;wire n5400_t;wire n5401;wire n5401_t;wire n5402;wire n5402_t;wire n5403;wire n5403_t;wire n5404;wire n5404_t;wire n5405;wire n5405_t;wire n5406;wire n5406_t;wire n5407;wire n5407_t;wire n5408;wire n5408_t;wire n5409;wire n5409_t;wire n5410;wire n5410_t;wire n5411;wire n5411_t;wire n5412;wire n5412_t;wire n5413;wire n5413_t;wire n5414;wire n5414_t;wire n5415;wire n5415_t;wire n5416;wire n5416_t;wire n5417;wire n5417_t;wire n5418;wire n5418_t;wire n5419;wire n5419_t;wire n5420;wire n5420_t;wire n5421;wire n5421_t;wire n5422;wire n5422_t;wire n5423;wire n5423_t;wire n5424;wire n5424_t;wire n5425;wire n5425_t;wire n5426;wire n5426_t;wire n5427;wire n5427_t;wire n5428;wire n5428_t;wire n5429;wire n5429_t;wire n5430;wire n5430_t;wire n5431;wire n5431_t;wire n5432;wire n5432_t;wire n5433;wire n5433_t;wire n5434;wire n5434_t;wire n5435;wire n5435_t;wire n5436;wire n5436_t;wire n5437;wire n5437_t;wire n5438;wire n5438_t;wire n5439;wire n5439_t;wire n5440;wire n5440_t;wire n5441;wire n5441_t;wire n5442;wire n5442_t;wire n5443;wire n5443_t;wire n5444;wire n5444_t;wire n5445;wire n5445_t;wire n5446;wire n5446_t;wire n5447;wire n5447_t;wire n5448;wire n5448_t;wire n5449;wire n5449_t;wire n5450;wire n5450_t;wire n5451;wire n5451_t;wire n5452;wire n5452_t;wire n5453;wire n5453_t;wire n5454;wire n5454_t;wire n5455;wire n5455_t;wire n5456;wire n5456_t;wire n5457;wire n5457_t;wire n5458;wire n5458_t;wire n5459;wire n5459_t;wire n5460;wire n5460_t;wire n5461;wire n5461_t;wire n5462;wire n5462_t;wire n5463;wire n5463_t;wire n5464;wire n5464_t;wire n5465;wire n5465_t;wire n5466;wire n5466_t;wire n5467;wire n5467_t;wire n5468;wire n5468_t;wire n5469;wire n5469_t;wire n5470;wire n5470_t;wire n5471;wire n5471_t;wire n5472;wire n5472_t;wire n5473;wire n5473_t;wire n5474;wire n5474_t;wire n5475;wire n5475_t;wire n5476;wire n5476_t;wire n5477;wire n5477_t;wire n5478;wire n5478_t;wire n5479;wire n5479_t;wire n5480;wire n5480_t;wire n5481;wire n5481_t;wire n5482;wire n5482_t;wire n5483;wire n5483_t;wire n5484;wire n5484_t;wire n5485;wire n5485_t;wire n5486;wire n5486_t;wire n5487;wire n5487_t;wire n5488;wire n5488_t;wire n5489;wire n5489_t;wire n5490;wire n5490_t;wire n5491;wire n5491_t;wire n5492;wire n5492_t;wire n5493;wire n5493_t;wire n5494;wire n5494_t;wire n5495;wire n5495_t;wire n5496;wire n5496_t;wire n5497;wire n5497_t;wire n5498;wire n5498_t;wire n5499;wire n5499_t;wire n5500;wire n5500_t;wire n5501;wire n5501_t;wire n5502;wire n5502_t;wire n5503;wire n5503_t;wire n5504;wire n5504_t;wire n5505;wire n5505_t;wire n5506;wire n5506_t;wire n5507;wire n5507_t;wire n5508;wire n5508_t;wire n5509;wire n5509_t;wire n5510;wire n5510_t;wire n5511;wire n5511_t;wire n5512;wire n5512_t;wire n5513;wire n5513_t;wire n5514;wire n5514_t;wire n5515;wire n5515_t;wire n5516;wire n5516_t;wire n5517;wire n5517_t;wire n5518;wire n5518_t;wire n5519;wire n5519_t;wire n5520;wire n5520_t;wire n5521;wire n5521_t;wire n5522;wire n5522_t;wire n5523;wire n5523_t;wire n5524;wire n5524_t;wire n5525;wire n5525_t;wire n5526;wire n5526_t;wire n5527;wire n5527_t;wire n5528;wire n5528_t;wire n5529;wire n5529_t;wire n5530;wire n5530_t;wire n5531;wire n5531_t;wire n5532;wire n5532_t;wire n5533;wire n5533_t;wire n5534;wire n5534_t;wire n5535;wire n5535_t;wire n5536;wire n5536_t;wire n5537;wire n5537_t;wire n5538;wire n5538_t;wire n5539;wire n5539_t;wire n5540;wire n5540_t;wire n5541;wire n5541_t;wire n5542;wire n5542_t;wire n5543;wire n5543_t;wire n5544;wire n5544_t;wire n5545;wire n5545_t;wire n5546;wire n5546_t;wire n5547;wire n5547_t;wire n5548;wire n5548_t;wire n5549;wire n5549_t;wire n5550;wire n5550_t;wire n5551;wire n5551_t;wire n5552;wire n5552_t;wire n5553;wire n5553_t;wire n5554;wire n5554_t;wire n5555;wire n5555_t;wire n5556;wire n5556_t;wire n5557;wire n5557_t;wire n5558;wire n5558_t;wire n5559;wire n5559_t;wire n5560;wire n5560_t;wire n5561;wire n5561_t;wire n5562;wire n5562_t;wire n5563;wire n5563_t;wire n5564;wire n5564_t;wire n5565;wire n5565_t;wire n5566;wire n5566_t;wire n5567;wire n5567_t;wire n5568;wire n5568_t;wire n5569;wire n5569_t;wire n5570;wire n5570_t;wire n5571;wire n5571_t;wire n5572;wire n5572_t;wire n5573;wire n5573_t;wire n5574;wire n5574_t;wire n5575;wire n5575_t;wire n5576;wire n5576_t;wire n5577;wire n5577_t;wire n5578;wire n5578_t;wire n5579;wire n5579_t;wire n5580;wire n5580_t;wire n5581;wire n5581_t;wire n5582;wire n5582_t;wire n5583;wire n5583_t;wire n5584;wire n5584_t;wire n5585;wire n5585_t;wire n5586;wire n5586_t;wire n5587;wire n5587_t;wire n5588;wire n5588_t;wire n5589;wire n5589_t;wire n5590;wire n5590_t;wire n5591;wire n5591_t;wire n5592;wire n5592_t;wire n5593;wire n5593_t;wire n5594;wire n5594_t;wire n5595;wire n5595_t;wire n5596;wire n5596_t;wire n5597;wire n5597_t;wire n5598;wire n5598_t;wire n5599;wire n5599_t;wire n5600;wire n5600_t;wire n5601;wire n5601_t;wire n5602;wire n5602_t;wire n5603;wire n5603_t;wire n5604;wire n5604_t;wire n5605;wire n5605_t;wire n5606;wire n5606_t;wire n5607;wire n5607_t;wire n5608;wire n5608_t;wire n5609;wire n5609_t;wire n5610;wire n5610_t;wire n5611;wire n5611_t;wire n5612;wire n5612_t;wire n5613;wire n5613_t;wire n5614;wire n5614_t;wire n5615;wire n5615_t;wire n5616;wire n5616_t;wire n5617;wire n5617_t;wire n5618;wire n5618_t;wire n5619;wire n5619_t;wire n5620;wire n5620_t;wire n5621;wire n5621_t;wire n5622;wire n5622_t;wire n5623;wire n5623_t;wire n5624;wire n5624_t;wire n5625;wire n5625_t;wire n5626;wire n5626_t;wire n5627;wire n5627_t;wire n5628;wire n5628_t;wire n5629;wire n5629_t;wire n5630;wire n5630_t;wire n5631;wire n5631_t;wire n5632;wire n5632_t;wire n5633;wire n5633_t;wire n5634;wire n5634_t;wire n5635;wire n5635_t;wire n5636;wire n5636_t;wire n5637;wire n5637_t;wire n5638;wire n5638_t;wire n5639;wire n5639_t;wire n5640;wire n5640_t;wire n5641;wire n5641_t;wire n5642;wire n5642_t;wire n5643;wire n5643_t;wire n5644;wire n5644_t;wire n5645;wire n5645_t;wire n5646;wire n5646_t;wire n5647;wire n5647_t;wire n5648;wire n5648_t;wire n5649;wire n5649_t;wire n5650;wire n5650_t;wire n5651;wire n5651_t;wire n5652;wire n5652_t;wire n5653;wire n5653_t;wire n5654;wire n5654_t;wire n5655;wire n5655_t;wire n5656;wire n5656_t;wire n5657;wire n5657_t;wire n5658;wire n5658_t;wire n5659;wire n5659_t;wire n5660;wire n5660_t;wire n5661;wire n5661_t;wire n5662;wire n5662_t;wire n5663;wire n5663_t;wire n5664;wire n5664_t;wire n5665;wire n5665_t;wire n5666;wire n5666_t;wire n5667;wire n5667_t;wire n5668;wire n5668_t;wire n5669;wire n5669_t;wire n5670;wire n5670_t;wire n5671;wire n5671_t;wire n5672;wire n5672_t;wire n5673;wire n5673_t;wire n5674;wire n5674_t;wire n5675;wire n5675_t;wire n5676;wire n5676_t;wire n5677;wire n5677_t;wire n5678;wire n5678_t;wire n5679;wire n5679_t;wire n5680;wire n5680_t;wire n5681;wire n5681_t;wire n5682;wire n5682_t;wire n5683;wire n5683_t;wire n5684;wire n5684_t;wire n5685;wire n5685_t;wire n5686;wire n5686_t;wire n5687;wire n5687_t;wire n5688;wire n5688_t;wire n5689;wire n5689_t;wire n5690;wire n5690_t;wire n5691;wire n5691_t;wire n5692;wire n5692_t;wire n5693;wire n5693_t;wire n5694;wire n5694_t;wire n5695;wire n5695_t;wire n5696;wire n5696_t;wire n5697;wire n5697_t;wire n5698;wire n5698_t;wire n5699;wire n5699_t;wire n5700;wire n5700_t;wire n5701;wire n5701_t;wire n5702;wire n5702_t;wire n5703;wire n5703_t;wire n5704;wire n5704_t;wire n5705;wire n5705_t;wire n5706;wire n5706_t;wire n5707;wire n5707_t;wire n5708;wire n5708_t;wire n5709;wire n5709_t;wire n5710;wire n5710_t;wire n5711;wire n5711_t;wire n5712;wire n5712_t;wire n5713;wire n5713_t;wire n5714;wire n5714_t;wire n5715;wire n5715_t;wire n5716;wire n5716_t;wire n5717;wire n5717_t;wire n5718;wire n5718_t;wire n5719;wire n5719_t;wire n5720;wire n5720_t;wire n5721;wire n5721_t;wire n5722;wire n5722_t;wire n5723;wire n5723_t;wire n5724;wire n5724_t;wire n5725;wire n5725_t;wire n5726;wire n5726_t;wire n5727;wire n5727_t;wire n5728;wire n5728_t;wire n5729;wire n5729_t;wire n5730;wire n5730_t;wire n5731;wire n5731_t;wire n5732;wire n5732_t;wire n5733;wire n5733_t;wire n5734;wire n5734_t;wire n5735;wire n5735_t;wire n5736;wire n5736_t;wire n5737;wire n5737_t;wire n5738;wire n5738_t;wire n5739;wire n5739_t;wire n5740;wire n5740_t;wire n5741;wire n5741_t;wire n5742;wire n5742_t;wire n5743;wire n5743_t;wire n5744;wire n5744_t;wire n5745;wire n5745_t;wire n5746;wire n5746_t;wire n5747;wire n5747_t;wire n5748;wire n5748_t;wire n5749;wire n5749_t;wire n5750;wire n5750_t;wire n5751;wire n5751_t;wire n5752;wire n5752_t;wire n5753;wire n5753_t;wire n5754;wire n5754_t;wire n5755;wire n5755_t;wire n5756;wire n5756_t;wire n5757;wire n5757_t;wire n5758;wire n5758_t;wire n5759;wire n5759_t;wire n5760;wire n5760_t;wire n5761;wire n5761_t;wire n5762;wire n5762_t;wire n5763;wire n5763_t;wire n5764;wire n5764_t;wire n5765;wire n5765_t;wire n5766;wire n5766_t;wire n5767;wire n5767_t;wire n5768;wire n5768_t;wire n5769;wire n5769_t;wire n5770;wire n5770_t;wire n5771;wire n5771_t;wire n5772;wire n5772_t;wire n5773;wire n5773_t;wire n5774;wire n5774_t;wire n5775;wire n5775_t;wire n5776;wire n5776_t;wire n5777;wire n5777_t;wire n5778;wire n5778_t;wire n5779;wire n5779_t;wire n5780;wire n5780_t;wire n5781;wire n5781_t;wire n5782;wire n5782_t;wire n5783;wire n5783_t;wire n5784;wire n5784_t;wire n5785;wire n5785_t;wire n5786;wire n5786_t;wire n5787;wire n5787_t;wire n5788;wire n5788_t;wire n5789;wire n5789_t;wire n5790;wire n5790_t;wire n5791;wire n5791_t;wire n5792;wire n5792_t;wire n5793;wire n5793_t;wire n5794;wire n5794_t;wire n5795;wire n5795_t;wire n5796;wire n5796_t;wire n5797;wire n5797_t;wire n5798;wire n5798_t;wire n5799;wire n5799_t;wire n5800;wire n5800_t;wire n5801;wire n5801_t;wire n5802;wire n5802_t;wire n5803;wire n5803_t;wire n5804;wire n5804_t;wire n5805;wire n5805_t;wire n5806;wire n5806_t;wire n5807;wire n5807_t;wire n5808;wire n5808_t;wire n5809;wire n5809_t;wire n5810;wire n5810_t;wire n5811;wire n5811_t;wire n5812;wire n5812_t;wire n5813;wire n5813_t;wire n5814;wire n5814_t;wire n5815;wire n5815_t;wire n5816;wire n5816_t;wire n5817;wire n5817_t;wire n5818;wire n5818_t;wire n5819;wire n5819_t;wire n5820;wire n5820_t;wire n5821;wire n5821_t;wire n5822;wire n5822_t;wire n5823;wire n5823_t;wire n5824;wire n5824_t;wire n5825;wire n5825_t;wire n5826;wire n5826_t;wire n5827;wire n5827_t;wire n5828;wire n5828_t;wire n5829;wire n5829_t;wire n5830;wire n5830_t;wire n5831;wire n5831_t;wire n5832;wire n5832_t;wire n5833;wire n5833_t;wire n5834;wire n5834_t;wire n5835;wire n5835_t;wire n5836;wire n5836_t;wire n5837;wire n5837_t;wire n5838;wire n5838_t;wire n5839;wire n5839_t;wire n5840;wire n5840_t;wire n5841;wire n5841_t;wire n5842;wire n5842_t;wire n5843;wire n5843_t;wire n5844;wire n5844_t;wire n5845;wire n5845_t;wire n5846;wire n5846_t;wire n5847;wire n5847_t;wire n5848;wire n5848_t;wire n5849;wire n5849_t;wire n5850;wire n5850_t;wire n5851;wire n5851_t;wire n5852;wire n5852_t;wire n5853;wire n5853_t;wire n5854;wire n5854_t;wire n5855;wire n5855_t;wire n5856;wire n5856_t;wire n5857;wire n5857_t;wire n5858;wire n5858_t;wire n5859;wire n5859_t;wire n5860;wire n5860_t;wire n5861;wire n5861_t;wire n5862;wire n5862_t;wire n5863;wire n5863_t;wire n5864;wire n5864_t;wire n5865;wire n5865_t;wire n5866;wire n5866_t;wire n5867;wire n5867_t;wire n5868;wire n5868_t;wire n5869;wire n5869_t;wire n5870;wire n5870_t;wire n5871;wire n5871_t;wire n5872;wire n5872_t;wire n5873;wire n5873_t;wire n5874;wire n5874_t;wire n5875;wire n5875_t;wire n5876;wire n5876_t;wire n5877;wire n5877_t;wire n5878;wire n5878_t;wire n5879;wire n5879_t;wire n5880;wire n5880_t;wire n5881;wire n5881_t;wire n5882;wire n5882_t;wire n5883;wire n5883_t;wire n5884;wire n5884_t;wire n5885;wire n5885_t;wire n5886;wire n5886_t;wire n5887;wire n5887_t;wire n5888;wire n5888_t;wire n5889;wire n5889_t;wire n5890;wire n5890_t;wire n5891;wire n5891_t;wire n5892;wire n5892_t;wire n5893;wire n5893_t;wire n5894;wire n5894_t;wire n5895;wire n5895_t;wire n5896;wire n5896_t;wire n5897;wire n5897_t;wire n5898;wire n5898_t;wire n5899;wire n5899_t;wire n5900;wire n5900_t;wire n5901;wire n5901_t;wire n5902;wire n5902_t;wire n5903;wire n5903_t;wire n5904;wire n5904_t;wire n5905;wire n5905_t;wire n5906;wire n5906_t;wire n5907;wire n5907_t;wire n5908;wire n5908_t;wire n5909;wire n5909_t;wire n5910;wire n5910_t;wire n5911;wire n5911_t;wire n5912;wire n5912_t;wire n5913;wire n5913_t;wire n5914;wire n5914_t;wire n5915;wire n5915_t;wire n5916;wire n5916_t;wire n5917;wire n5917_t;wire n5918;wire n5918_t;wire n5919;wire n5919_t;wire n5920;wire n5920_t;wire n5921;wire n5921_t;wire n5922;wire n5922_t;wire n5923;wire n5923_t;wire n5924;wire n5924_t;wire n5925;wire n5925_t;wire n5926;wire n5926_t;wire n5927;wire n5927_t;wire n5928;wire n5928_t;wire n5929;wire n5929_t;wire n5930;wire n5930_t;wire n5931;wire n5931_t;wire n5932;wire n5932_t;wire n5933;wire n5933_t;wire n5934;wire n5934_t;wire n5935;wire n5935_t;wire n5936;wire n5936_t;wire n5937;wire n5937_t;wire n5938;wire n5938_t;wire n5939;wire n5939_t;wire n5940;wire n5940_t;wire n5941;wire n5941_t;wire n5942;wire n5942_t;wire n5943;wire n5943_t;wire n5944;wire n5944_t;wire n5945;wire n5945_t;wire n5946;wire n5946_t;wire n5947;wire n5947_t;wire n5948;wire n5948_t;wire n5949;wire n5949_t;wire n5950;wire n5950_t;wire n5951;wire n5951_t;wire n5952;wire n5952_t;wire n5953;wire n5953_t;wire n5954;wire n5954_t;wire n5955;wire n5955_t;wire n5956;wire n5956_t;wire n5957;wire n5957_t;wire n5958;wire n5958_t;wire n5959;wire n5959_t;wire n5960;wire n5960_t;wire n5961;wire n5961_t;wire n5962;wire n5962_t;wire n5963;wire n5963_t;wire n5964;wire n5964_t;wire n5965;wire n5965_t;wire n5966;wire n5966_t;wire n5967;wire n5967_t;wire n5968;wire n5968_t;wire n5969;wire n5969_t;wire n5970;wire n5970_t;wire n5971;wire n5971_t;wire n5972;wire n5972_t;wire n5973;wire n5973_t;wire n5974;wire n5974_t;wire n5975;wire n5975_t;wire n5976;wire n5976_t;wire n5977;wire n5977_t;wire n5978;wire n5978_t;wire n5979;wire n5979_t;wire n5980;wire n5980_t;wire n5981;wire n5981_t;wire n5982;wire n5982_t;wire n5983;wire n5983_t;wire n5984;wire n5984_t;wire n5985;wire n5985_t;wire n5986;wire n5986_t;wire n5987;wire n5987_t;wire n5988;wire n5988_t;wire n5989;wire n5989_t;wire n5990;wire n5990_t;wire n5991;wire n5991_t;wire n5992;wire n5992_t;wire n5993;wire n5993_t;wire n5994;wire n5994_t;wire n5995;wire n5995_t;wire n5996;wire n5996_t;wire n5997;wire n5997_t;wire n5998;wire n5998_t;wire n5999;wire n5999_t;wire n6000;wire n6000_t;wire n6001;wire n6001_t;wire n6002;wire n6002_t;wire n6003;wire n6003_t;wire n6004;wire n6004_t;wire n6005;wire n6005_t;wire n6006;wire n6006_t;wire n6007;wire n6007_t;wire n6008;wire n6008_t;wire n6009;wire n6009_t;wire n6010;wire n6010_t;wire n6011;wire n6011_t;wire n6012;wire n6012_t;wire n6013;wire n6013_t;wire n6014;wire n6014_t;wire n6015;wire n6015_t;wire n6016;wire n6016_t;wire n6017;wire n6017_t;wire n6018;wire n6018_t;wire n6019;wire n6019_t;wire n6020;wire n6020_t;wire n6021;wire n6021_t;wire n6022;wire n6022_t;wire n6023;wire n6023_t;wire n6024;wire n6024_t;wire n6025;wire n6025_t;wire n6026;wire n6026_t;wire n6027;wire n6027_t;wire n6028;wire n6028_t;wire n6029;wire n6029_t;wire n6030;wire n6030_t;wire n6031;wire n6031_t;wire n6032;wire n6032_t;wire n6033;wire n6033_t;wire n6034;wire n6034_t;wire n6035;wire n6035_t;wire n6036;wire n6036_t;wire n6037;wire n6037_t;wire n6038;wire n6038_t;wire n6039;wire n6039_t;wire n6040;wire n6040_t;wire n6041;wire n6041_t;wire n6042;wire n6042_t;wire n6043;wire n6043_t;wire n6044;wire n6044_t;wire n6045;wire n6045_t;wire n6046;wire n6046_t;wire n6047;wire n6047_t;wire n6048;wire n6048_t;wire n6049;wire n6049_t;wire n6050;wire n6050_t;wire n6051;wire n6051_t;wire n6052;wire n6052_t;wire n6053;wire n6053_t;wire n6054;wire n6054_t;wire n6055;wire n6055_t;wire n6056;wire n6056_t;wire n6057;wire n6057_t;wire n6058;wire n6058_t;wire n6059;wire n6059_t;wire n6060;wire n6060_t;wire n6061;wire n6061_t;wire n6062;wire n6062_t;wire n6063;wire n6063_t;wire n6064;wire n6064_t;wire n6065;wire n6065_t;wire n6066;wire n6066_t;wire n6067;wire n6067_t;wire n6068;wire n6068_t;wire n6069;wire n6069_t;wire n6070;wire n6070_t;wire n6071;wire n6071_t;wire n6072;wire n6072_t;wire n6073;wire n6073_t;wire n6074;wire n6074_t;wire n6075;wire n6075_t;wire n6076;wire n6076_t;wire n6077;wire n6077_t;wire n6078;wire n6078_t;wire n6079;wire n6079_t;wire n6080;wire n6080_t;wire n6081;wire n6081_t;wire n6082;wire n6082_t;wire n6083;wire n6083_t;wire n6084;wire n6084_t;wire n6085;wire n6085_t;wire n6086;wire n6086_t;wire n6087;wire n6087_t;wire n6088;wire n6088_t;wire n6089;wire n6089_t;wire n6090;wire n6090_t;wire n6091;wire n6091_t;wire n6092;wire n6092_t;wire n6093;wire n6093_t;wire n6094;wire n6094_t;wire n6095;wire n6095_t;wire n6096;wire n6096_t;wire n6097;wire n6097_t;wire n6098;wire n6098_t;wire n6099;wire n6099_t;wire n6100;wire n6100_t;wire n6101;wire n6101_t;wire n6102;wire n6102_t;wire n6103;wire n6103_t;wire n6104;wire n6104_t;wire n6105;wire n6105_t;wire n6106;wire n6106_t;wire n6107;wire n6107_t;wire n6108;wire n6108_t;wire n6109;wire n6109_t;wire n6110;wire n6110_t;wire n6111;wire n6111_t;wire n6112;wire n6112_t;wire n6113;wire n6113_t;wire n6114;wire n6114_t;wire n6115;wire n6115_t;wire n6116;wire n6116_t;wire n6117;wire n6117_t;wire n6118;wire n6118_t;wire n6119;wire n6119_t;wire n6120;wire n6120_t;wire n6121;wire n6121_t;wire n6122;wire n6122_t;wire n6123;wire n6123_t;wire n6124;wire n6124_t;wire n6125;wire n6125_t;wire n6126;wire n6126_t;wire n6127;wire n6127_t;wire n6128;wire n6128_t;wire n6129;wire n6129_t;wire n6130;wire n6130_t;wire n6131;wire n6131_t;wire n6132;wire n6132_t;wire n6133;wire n6133_t;wire n6134;wire n6134_t;wire n6135;wire n6135_t;wire n6136;wire n6136_t;wire n6137;wire n6137_t;wire n6138;wire n6138_t;wire n6139;wire n6139_t;wire n6140;wire n6140_t;wire n6141;wire n6141_t;wire n6142;wire n6142_t;wire n6143;wire n6143_t;wire n6144;wire n6144_t;wire n6145;wire n6145_t;wire n6146;wire n6146_t;wire n6147;wire n6147_t;wire n6148;wire n6148_t;wire n6149;wire n6149_t;wire n6150;wire n6150_t;wire n6151;wire n6151_t;wire n6152;wire n6152_t;wire n6153;wire n6153_t;wire n6154;wire n6154_t;wire n6155;wire n6155_t;wire n6156;wire n6156_t;wire n6157;wire n6157_t;wire n6158;wire n6158_t;wire n6159;wire n6159_t;wire n6160;wire n6160_t;wire n6161;wire n6161_t;wire n6162;wire n6162_t;wire n6163;wire n6163_t;wire n6164;wire n6164_t;wire n6165;wire n6165_t;wire n6166;wire n6166_t;wire n6167;wire n6167_t;wire n6168;wire n6168_t;wire n6169;wire n6169_t;wire n6170;wire n6170_t;wire n6171;wire n6171_t;wire n6172;wire n6172_t;wire n6173;wire n6173_t;wire n6174;wire n6174_t;wire n6175;wire n6175_t;wire n6176;wire n6176_t;wire n6177;wire n6177_t;wire n6178;wire n6178_t;wire n6179;wire n6179_t;wire n6180;wire n6180_t;wire n6181;wire n6181_t;wire n6182;wire n6182_t;wire n6183;wire n6183_t;wire n6184;wire n6184_t;wire n6185;wire n6185_t;wire n6186;wire n6186_t;wire n6187;wire n6187_t;wire n6188;wire n6188_t;wire n6189;wire n6189_t;wire n6190;wire n6190_t;wire n6191;wire n6191_t;wire n6192;wire n6192_t;wire n6193;wire n6193_t;wire n6194;wire n6194_t;wire n6195;wire n6195_t;wire n6196;wire n6196_t;wire n6197;wire n6197_t;wire n6198;wire n6198_t;wire n6199;wire n6199_t;wire n6200;wire n6200_t;wire n6201;wire n6201_t;wire n6202;wire n6202_t;wire n6203;wire n6203_t;wire n6204;wire n6204_t;wire n6205;wire n6205_t;wire n6206;wire n6206_t;wire n6207;wire n6207_t;wire n6208;wire n6208_t;wire n6209;wire n6209_t;wire n6210;wire n6210_t;wire n6211;wire n6211_t;wire n6212;wire n6212_t;wire n6213;wire n6213_t;wire n6214;wire n6214_t;wire n6215;wire n6215_t;wire n6216;wire n6216_t;wire n6217;wire n6217_t;wire n6218;wire n6218_t;wire n6219;wire n6219_t;wire n6220;wire n6220_t;wire n6221;wire n6221_t;wire n6222;wire n6222_t;wire n6223;wire n6223_t;wire n6224;wire n6224_t;wire n6225;wire n6225_t;wire n6226;wire n6226_t;wire n6227;wire n6227_t;wire n6228;wire n6228_t;wire n6229;wire n6229_t;wire n6230;wire n6230_t;wire n6231;wire n6231_t;wire n6232;wire n6232_t;wire n6233;wire n6233_t;wire n6234;wire n6234_t;wire n6235;wire n6235_t;wire n6236;wire n6236_t;wire n6237;wire n6237_t;wire n6238;wire n6238_t;wire n6239;wire n6239_t;wire n6240;wire n6240_t;wire n6241;wire n6241_t;wire n6242;wire n6242_t;wire n6243;wire n6243_t;wire n6244;wire n6244_t;wire n6245;wire n6245_t;wire n6246;wire n6246_t;wire n6247;wire n6247_t;wire n6248;wire n6248_t;wire n6249;wire n6249_t;wire n6250;wire n6250_t;wire n6251;wire n6251_t;wire n6252;wire n6252_t;wire n6253;wire n6253_t;wire n6254;wire n6254_t;wire n6255;wire n6255_t;wire n6256;wire n6256_t;wire n6257;wire n6257_t;wire n6258;wire n6258_t;wire n6259;wire n6259_t;wire n6260;wire n6260_t;wire n6261;wire n6261_t;wire n6262;wire n6262_t;wire n6263;wire n6263_t;wire n6264;wire n6264_t;wire n6265;wire n6265_t;wire n6266;wire n6266_t;wire n6267;wire n6267_t;wire n6268;wire n6268_t;wire n6269;wire n6269_t;wire n6270;wire n6270_t;wire n6271;wire n6271_t;wire n6272;wire n6272_t;wire n6273;wire n6273_t;wire n6274;wire n6274_t;wire n6275;wire n6275_t;wire n6276;wire n6276_t;wire n6277;wire n6277_t;wire n6278;wire n6278_t;wire n6279;wire n6279_t;wire n6280;wire n6280_t;wire n6281;wire n6281_t;wire n6282;wire n6282_t;wire n6283;wire n6283_t;wire n6284;wire n6284_t;wire n6285;wire n6285_t;wire n6286;wire n6286_t;wire n6287;wire n6287_t;wire n6288;wire n6288_t;wire n6289;wire n6289_t;wire n6290;wire n6290_t;wire n6291;wire n6291_t;wire n6292;wire n6292_t;wire n6293;wire n6293_t;wire n6294;wire n6294_t;wire n6295;wire n6295_t;wire n6296;wire n6296_t;wire n6297;wire n6297_t;wire n6298;wire n6298_t;wire n6299;wire n6299_t;wire n6300;wire n6300_t;wire n6301;wire n6301_t;wire n6302;wire n6302_t;wire n6303;wire n6303_t;wire n6304;wire n6304_t;wire n6305;wire n6305_t;wire n6306;wire n6306_t;wire n6307;wire n6307_t;wire n6308;wire n6308_t;wire n6309;wire n6309_t;wire n6310;wire n6310_t;wire n6311;wire n6311_t;wire n6312;wire n6312_t;wire n6313;wire n6313_t;wire n6314;wire n6314_t;wire n6315;wire n6315_t;wire n6316;wire n6316_t;wire n6317;wire n6317_t;wire n6318;wire n6318_t;wire n6319;wire n6319_t;wire n6320;wire n6320_t;wire n6321;wire n6321_t;wire n6322;wire n6322_t;wire n6323;wire n6323_t;wire n6324;wire n6324_t;wire n6325;wire n6325_t;wire n6326;wire n6326_t;wire n6327;wire n6327_t;wire n6328;wire n6328_t;wire n6329;wire n6329_t;wire n6330;wire n6330_t;wire n6331;wire n6331_t;wire n6332;wire n6332_t;wire n6333;wire n6333_t;wire n6334;wire n6334_t;wire n6335;wire n6335_t;wire n6336;wire n6336_t;wire n6337;wire n6337_t;wire n6338;wire n6338_t;wire n6339;wire n6339_t;wire n6340;wire n6340_t;wire n6341;wire n6341_t;wire n6342;wire n6342_t;wire n6343;wire n6343_t;wire n6344;wire n6344_t;wire n6345;wire n6345_t;wire n6346;wire n6346_t;wire n6347;wire n6347_t;wire n6348;wire n6348_t;wire n6349;wire n6349_t;wire n6350;wire n6350_t;wire n6351;wire n6351_t;wire n6352;wire n6352_t;wire n6353;wire n6353_t;wire n6354;wire n6354_t;wire n6355;wire n6355_t;wire n6356;wire n6356_t;wire n6357;wire n6357_t;wire n6358;wire n6358_t;wire n6359;wire n6359_t;wire n6360;wire n6360_t;wire n6361;wire n6361_t;wire n6362;wire n6362_t;wire n6363;wire n6363_t;wire n6364;wire n6364_t;wire n6365;wire n6365_t;wire n6366;wire n6366_t;wire n6367;wire n6367_t;wire n6368;wire n6368_t;wire n6369;wire n6369_t;wire n6370;wire n6370_t;wire n6371;wire n6371_t;wire n6372;wire n6372_t;wire n6373;wire n6373_t;wire n6374;wire n6374_t;wire n6375;wire n6375_t;wire n6376;wire n6376_t;wire n6377;wire n6377_t;wire n6378;wire n6378_t;wire n6379;wire n6379_t;wire n6380;wire n6380_t;wire n6381;wire n6381_t;wire n6382;wire n6382_t;wire n6383;wire n6383_t;wire n6384;wire n6384_t;wire n6385;wire n6385_t;wire n6386;wire n6386_t;wire n6387;wire n6387_t;wire n6388;wire n6388_t;wire n6389;wire n6389_t;wire n6390;wire n6390_t;wire n6391;wire n6391_t;wire n6392;wire n6392_t;wire n6393;wire n6393_t;wire n6394;wire n6394_t;wire n6395;wire n6395_t;wire n6396;wire n6396_t;wire n6397;wire n6397_t;wire n6398;wire n6398_t;wire n6399;wire n6399_t;wire n6400;wire n6400_t;wire n6401;wire n6401_t;wire n6402;wire n6402_t;wire n6403;wire n6403_t;wire n6404;wire n6404_t;wire n6405;wire n6405_t;wire n6406;wire n6406_t;wire n6407;wire n6407_t;wire n6408;wire n6408_t;wire n6409;wire n6409_t;wire n6410;wire n6410_t;wire n6411;wire n6411_t;wire n6412;wire n6412_t;wire n6413;wire n6413_t;wire n6414;wire n6414_t;wire n6415;wire n6415_t;wire n6416;wire n6416_t;wire n6417;wire n6417_t;wire n6418;wire n6418_t;wire n6419;wire n6419_t;wire n6420;wire n6420_t;wire n6421;wire n6421_t;wire n6422;wire n6422_t;wire n6423;wire n6423_t;wire n6424;wire n6424_t;wire n6425;wire n6425_t;wire n6426;wire n6426_t;wire n6427;wire n6427_t;wire n6428;wire n6428_t;wire n6429;wire n6429_t;wire n6430;wire n6430_t;wire n6431;wire n6431_t;wire n6432;wire n6432_t;wire n6433;wire n6433_t;wire n6434;wire n6434_t;wire n6435;wire n6435_t;wire n6436;wire n6436_t;wire n6437;wire n6437_t;wire n6438;wire n6438_t;wire n6439;wire n6439_t;wire n6440;wire n6440_t;wire n6441;wire n6441_t;wire n6442;wire n6442_t;wire n6443;wire n6443_t;wire n6444;wire n6444_t;wire n6445;wire n6445_t;wire n6446;wire n6446_t;wire n6447;wire n6447_t;wire n6448;wire n6448_t;wire n6449;wire n6449_t;wire n6450;wire n6450_t;wire n6451;wire n6451_t;wire n6452;wire n6452_t;wire n6453;wire n6453_t;wire n6454;wire n6454_t;wire n6455;wire n6455_t;wire n6456;wire n6456_t;wire n6457;wire n6457_t;wire n6458;wire n6458_t;wire n6459;wire n6459_t;wire n6460;wire n6460_t;wire n6461;wire n6461_t;wire n6462;wire n6462_t;wire n6463;wire n6463_t;wire n6464;wire n6464_t;wire n6465;wire n6465_t;wire n6466;wire n6466_t;wire n6467;wire n6467_t;wire n6468;wire n6468_t;wire n6469;wire n6469_t;wire n6470;wire n6470_t;wire n6471;wire n6471_t;wire n6472;wire n6472_t;wire n6473;wire n6473_t;wire n6474;wire n6474_t;wire n6475;wire n6475_t;wire n6476;wire n6476_t;wire n6477;wire n6477_t;wire n6478;wire n6478_t;wire n6479;wire n6479_t;wire n6480;wire n6480_t;wire n6481;wire n6481_t;wire n6482;wire n6482_t;wire n6483;wire n6483_t;wire n6484;wire n6484_t;wire n6485;wire n6485_t;wire n6486;wire n6486_t;wire n6487;wire n6487_t;wire n6488;wire n6488_t;wire n6489;wire n6489_t;wire n6490;wire n6490_t;wire n6491;wire n6491_t;wire n6492;wire n6492_t;wire n6493;wire n6493_t;wire n6494;wire n6494_t;wire n6495;wire n6495_t;wire n6496;wire n6496_t;wire n6497;wire n6497_t;wire n6498;wire n6498_t;wire n6499;wire n6499_t;wire n6500;wire n6500_t;wire n6501;wire n6501_t;wire n6502;wire n6502_t;wire n6503;wire n6503_t;wire n6504;wire n6504_t;wire n6505;wire n6505_t;wire n6506;wire n6506_t;wire n6507;wire n6507_t;wire n6508;wire n6508_t;wire n6509;wire n6509_t;wire n6510;wire n6510_t;wire n6511;wire n6511_t;wire n6512;wire n6512_t;wire n6513;wire n6513_t;wire n6514;wire n6514_t;wire n6515;wire n6515_t;wire n6516;wire n6516_t;wire n6517;wire n6517_t;wire n6518;wire n6518_t;wire n6519;wire n6519_t;wire n6520;wire n6520_t;wire n6521;wire n6521_t;wire n6522;wire n6522_t;wire n6523;wire n6523_t;wire n6524;wire n6524_t;wire n6525;wire n6525_t;wire n6526;wire n6526_t;wire n6527;wire n6527_t;wire n6528;wire n6528_t;wire n6529;wire n6529_t;wire n6530;wire n6530_t;wire n6531;wire n6531_t;wire n6532;wire n6532_t;wire n6533;wire n6533_t;wire n6534;wire n6534_t;wire n6535;wire n6535_t;wire n6536;wire n6536_t;wire n6537;wire n6537_t;wire n6538;wire n6538_t;wire n6539;wire n6539_t;wire n6540;wire n6540_t;wire n6541;wire n6541_t;wire n6542;wire n6542_t;wire n6543;wire n6543_t;wire n6544;wire n6544_t;wire n6545;wire n6545_t;wire n6546;wire n6546_t;wire n6547;wire n6547_t;wire n6548;wire n6548_t;wire n6549;wire n6549_t;wire n6550;wire n6550_t;wire n6551;wire n6551_t;wire n6552;wire n6552_t;wire n6553;wire n6553_t;wire n6554;wire n6554_t;wire n6555;wire n6555_t;wire n6556;wire n6556_t;wire n6557;wire n6557_t;wire n6558;wire n6558_t;wire n6559;wire n6559_t;wire n6560;wire n6560_t;wire n6561;wire n6561_t;wire n6562;wire n6562_t;wire n6563;wire n6563_t;wire n6564;wire n6564_t;wire n6565;wire n6565_t;wire n6566;wire n6566_t;wire n6567;wire n6567_t;wire n6568;wire n6568_t;wire n6569;wire n6569_t;wire n6570;wire n6570_t;wire n6571;wire n6571_t;wire n6572;wire n6572_t;wire n6573;wire n6573_t;wire n6574;wire n6574_t;wire n6575;wire n6575_t;wire n6576;wire n6576_t;wire n6577;wire n6577_t;wire n6578;wire n6578_t;wire n6579;wire n6579_t;wire n6580;wire n6580_t;wire n6581;wire n6581_t;wire n6582;wire n6582_t;wire n6583;wire n6583_t;wire n6584;wire n6584_t;wire n6585;wire n6585_t;wire n6586;wire n6586_t;wire n6587;wire n6587_t;wire n6588;wire n6588_t;wire n6589;wire n6589_t;wire n6590;wire n6590_t;wire n6591;wire n6591_t;wire n6592;wire n6592_t;wire n6593;wire n6593_t;wire n6594;wire n6594_t;wire n6595;wire n6595_t;wire n6596;wire n6596_t;wire n6597;wire n6597_t;wire n6598;wire n6598_t;wire n6599;wire n6599_t;wire n6600;wire n6600_t;wire n6601;wire n6601_t;wire n6602;wire n6602_t;wire n6603;wire n6603_t;wire n6604;wire n6604_t;wire n6605;wire n6605_t;wire n6606;wire n6606_t;wire n6607;wire n6607_t;wire n6608;wire n6608_t;wire n6609;wire n6609_t;wire n6610;wire n6610_t;wire n6611;wire n6611_t;wire n6612;wire n6612_t;wire n6613;wire n6613_t;wire n6614;wire n6614_t;wire n6615;wire n6615_t;wire n6616;wire n6616_t;wire n6617;wire n6617_t;wire n6618;wire n6618_t;wire n6619;wire n6619_t;wire n6620;wire n6620_t;wire n6621;wire n6621_t;wire n6622;wire n6622_t;wire n6623;wire n6623_t;wire n6624;wire n6624_t;wire n6625;wire n6625_t;wire n6626;wire n6626_t;wire n6627;wire n6627_t;wire n6628;wire n6628_t;wire n6629;wire n6629_t;wire n6630;wire n6630_t;wire n6631;wire n6631_t;wire n6632;wire n6632_t;wire n6633;wire n6633_t;wire n6634;wire n6634_t;wire n6635;wire n6635_t;wire n6636;wire n6636_t;wire n6637;wire n6637_t;wire n6638;wire n6638_t;wire n6639;wire n6639_t;wire n6640;wire n6640_t;wire n6641;wire n6641_t;wire n6642;wire n6642_t;wire n6643;wire n6643_t;wire n6644;wire n6644_t;wire n6645;wire n6645_t;wire n6646;wire n6646_t;wire n6647;wire n6647_t;wire n6648;wire n6648_t;wire n6649;wire n6649_t;wire n6650;wire n6650_t;wire n6651;wire n6651_t;wire n6652;wire n6652_t;wire n6653;wire n6653_t;wire n6654;wire n6654_t;wire n6655;wire n6655_t;wire n6656;wire n6656_t;wire n6657;wire n6657_t;wire n6658;wire n6658_t;wire n6659;wire n6659_t;wire n6660;wire n6660_t;wire n6661;wire n6661_t;wire n6662;wire n6662_t;wire n6663;wire n6663_t;wire n6664;wire n6664_t;wire n6665;wire n6665_t;wire n6666;wire n6666_t;wire n6667;wire n6667_t;wire n6668;wire n6668_t;wire n6669;wire n6669_t;wire n6670;wire n6670_t;wire n6671;wire n6671_t;wire n6672;wire n6672_t;wire n6673;wire n6673_t;wire n6674;wire n6674_t;wire n6675;wire n6675_t;wire n6676;wire n6676_t;wire n6677;wire n6677_t;wire n6678;wire n6678_t;wire n6679;wire n6679_t;wire n6680;wire n6680_t;wire n6681;wire n6681_t;wire n6682;wire n6682_t;wire n6683;wire n6683_t;wire n6684;wire n6684_t;wire n6685;wire n6685_t;wire n6686;wire n6686_t;wire n6687;wire n6687_t;wire n6688;wire n6688_t;wire n6689;wire n6689_t;wire n6690;wire n6690_t;wire n6691;wire n6691_t;wire n6692;wire n6692_t;wire n6693;wire n6693_t;wire n6694;wire n6694_t;wire n6695;wire n6695_t;wire n6696;wire n6696_t;wire n6697;wire n6697_t;wire n6698;wire n6698_t;wire n6699;wire n6699_t;wire n6700;wire n6700_t;wire n6701;wire n6701_t;wire n6702;wire n6702_t;wire n6703;wire n6703_t;wire n6704;wire n6704_t;wire n6705;wire n6705_t;wire n6706;wire n6706_t;wire n6707;wire n6707_t;wire n6708;wire n6708_t;wire n6709;wire n6709_t;wire n6710;wire n6710_t;wire n6711;wire n6711_t;wire n6712;wire n6712_t;wire n6713;wire n6713_t;wire n6714;wire n6714_t;wire n6715;wire n6715_t;wire n6716;wire n6716_t;wire n6717;wire n6717_t;wire n6718;wire n6718_t;wire n6719;wire n6719_t;wire n6720;wire n6720_t;wire n6721;wire n6721_t;wire n6722;wire n6722_t;wire n6723;wire n6723_t;wire n6724;wire n6724_t;wire n6725;wire n6725_t;wire n6726;wire n6726_t;wire n6727;wire n6727_t;wire n6728;wire n6728_t;wire n6729;wire n6729_t;wire n6730;wire n6730_t;wire n6731;wire n6731_t;wire n6732;wire n6732_t;wire n6733;wire n6733_t;wire n6734;wire n6734_t;wire n6735;wire n6735_t;wire n6736;wire n6736_t;wire n6737;wire n6737_t;wire n6738;wire n6738_t;wire n6739;wire n6739_t;wire n6740;wire n6740_t;wire n6741;wire n6741_t;wire n6742;wire n6742_t;wire n6743;wire n6743_t;wire n6744;wire n6744_t;wire n6745;wire n6745_t;wire n6746;wire n6746_t;wire n6747;wire n6747_t;wire n6748;wire n6748_t;wire n6749;wire n6749_t;wire n6750;wire n6750_t;wire n6751;wire n6751_t;wire n6752;wire n6752_t;wire n6753;wire n6753_t;wire n6754;wire n6754_t;wire n6755;wire n6755_t;wire n6756;wire n6756_t;wire n6757;wire n6757_t;wire n6758;wire n6758_t;wire n6759;wire n6759_t;wire n6760;wire n6760_t;wire n6761;wire n6761_t;wire n6762;wire n6762_t;wire n6763;wire n6763_t;wire n6764;wire n6764_t;wire n6765;wire n6765_t;wire n6766;wire n6766_t;wire n6767;wire n6767_t;wire n6768;wire n6768_t;wire n6769;wire n6769_t;wire n6770;wire n6770_t;wire n6771;wire n6771_t;wire n6772;wire n6772_t;wire n6773;wire n6773_t;wire n6774;wire n6774_t;wire n6775;wire n6775_t;wire n6776;wire n6776_t;wire n6777;wire n6777_t;wire n6778;wire n6778_t;wire n6779;wire n6779_t;wire n6780;wire n6780_t;wire n6781;wire n6781_t;wire n6782;wire n6782_t;wire n6783;wire n6783_t;wire n6784;wire n6784_t;wire n6785;wire n6785_t;wire n6786;wire n6786_t;wire n6787;wire n6787_t;wire n6788;wire n6788_t;wire n6789;wire n6789_t;wire n6790;wire n6790_t;wire n6791;wire n6791_t;wire n6792;wire n6792_t;wire n6793;wire n6793_t;wire n6794;wire n6794_t;wire n6795;wire n6795_t;wire n6796;wire n6796_t;wire n6797;wire n6797_t;wire n6798;wire n6798_t;wire n6799;wire n6799_t;wire n6800;wire n6800_t;wire n6801;wire n6801_t;wire n6802;wire n6802_t;wire n6803;wire n6803_t;wire n6804;wire n6804_t;wire n6805;wire n6805_t;wire n6806;wire n6806_t;wire n6807;wire n6807_t;wire n6808;wire n6808_t;wire n6811;wire n6811_t;wire n6812;wire n6812_t;wire n6813;wire n6813_t;wire n6814;wire n6814_t;wire n6815;wire n6815_t;wire n6816;wire n6816_t;wire n6817;wire n6817_t;wire n6818;wire n6818_t;wire n6819;wire n6819_t;wire n6820;wire n6820_t;wire n6821;wire n6821_t;wire n6822;wire n6822_t;wire n6823;wire n6823_t;wire n6824;wire n6824_t;wire n6825;wire n6825_t;wire n6826;wire n6826_t;wire n6827;wire n6827_t;wire n6828;wire n6828_t;wire n6829;wire n6829_t;wire n6830;wire n6830_t;wire n6831;wire n6831_t;wire n6832;wire n6832_t;wire n6833;wire n6833_t;wire n6834;wire n6834_t;wire n6835;wire n6835_t;wire n6836;wire n6836_t;wire n6837;wire n6837_t;wire n6838;wire n6838_t;wire n6839;wire n6839_t;wire n6840;wire n6840_t;wire n6841;wire n6841_t;wire n6842;wire n6842_t;wire n6843;wire n6843_t;wire n6844;wire n6844_t;wire n6845;wire n6845_t;wire n6846;wire n6846_t;wire n6847;wire n6847_t;wire n6848;wire n6848_t;wire n6849;wire n6849_t;wire n6850;wire n6850_t;wire n6851;wire n6851_t;wire n6852;wire n6852_t;wire n6853;wire n6853_t;wire n6854;wire n6854_t;wire n6855;wire n6855_t;wire n6856;wire n6856_t;wire n6857;wire n6857_t;wire n6858;wire n6858_t;wire n6859;wire n6859_t;wire n6860;wire n6860_t;wire n6861;wire n6861_t;wire n6862;wire n6862_t;wire n6863;wire n6863_t;wire n6864;wire n6864_t;wire n6865;wire n6865_t;wire n6866;wire n6866_t;wire n6867;wire n6867_t;wire n6868;wire n6868_t;wire n6869;wire n6869_t;wire n6870;wire n6870_t;wire n6871;wire n6871_t;wire n6872;wire n6872_t;wire n6873;wire n6873_t;wire n6874;wire n6874_t;wire n6875;wire n6875_t;wire n6876;wire n6876_t;wire n6877;wire n6877_t;wire n6878;wire n6878_t;wire n6879;wire n6879_t;wire n6880;wire n6880_t;wire n6881;wire n6881_t;wire n6882;wire n6882_t;wire n6883;wire n6883_t;wire n6884;wire n6884_t;wire n6885;wire n6885_t;wire n6886;wire n6886_t;wire n6887;wire n6887_t;wire n6888;wire n6888_t;wire n6889;wire n6889_t;wire n6890;wire n6890_t;wire n6891;wire n6891_t;wire n6892;wire n6892_t;wire n6893;wire n6893_t;wire n6894;wire n6894_t;wire n6895;wire n6895_t;wire n6896;wire n6896_t;wire n6897;wire n6897_t;wire n6898;wire n6898_t;wire n6899;wire n6899_t;wire n6900;wire n6900_t;wire n6901;wire n6901_t;wire n6902;wire n6902_t;wire n6903;wire n6903_t;wire n6904;wire n6904_t;wire n6905;wire n6905_t;wire n6906;wire n6906_t;wire n6907;wire n6907_t;wire n6908;wire n6908_t;wire n6909;wire n6909_t;wire n6910;wire n6910_t;wire n6911;wire n6911_t;wire n6912;wire n6912_t;wire n6913;wire n6913_t;wire n6914;wire n6914_t;wire n6915;wire n6915_t;wire n6916;wire n6916_t;wire n6917;wire n6917_t;wire n6918;wire n6918_t;wire n6919;wire n6919_t;wire n6920;wire n6920_t;wire n6921;wire n6921_t;wire n6922;wire n6922_t;wire n6923;wire n6923_t;wire n6924;wire n6924_t;wire n6925;wire n6925_t;wire n6926;wire n6926_t;wire n6927;wire n6927_t;wire n6928;wire n6928_t;wire n6929;wire n6929_t;wire n6930;wire n6930_t;wire n6931;wire n6931_t;wire n6932;wire n6932_t;wire n6933;wire n6933_t;wire n6934;wire n6934_t;wire n6935;wire n6935_t;wire n6936;wire n6936_t;wire n6937;wire n6937_t;wire n6938;wire n6938_t;wire n6939;wire n6939_t;wire n6940;wire n6940_t;wire n6941;wire n6941_t;wire n6942;wire n6942_t;wire n6943;wire n6943_t;wire n6944;wire n6944_t;wire n6945;wire n6945_t;wire n6946;wire n6946_t;wire n6947;wire n6947_t;wire n6948;wire n6948_t;wire n6949;wire n6949_t;wire n6950;wire n6950_t;wire n6951;wire n6951_t;wire n6952;wire n6952_t;wire n6953;wire n6953_t;wire n6954;wire n6954_t;wire n6955;wire n6955_t;wire n6956;wire n6956_t;wire n6957;wire n6957_t;wire n6958;wire n6958_t;wire n6959;wire n6959_t;wire n6960;wire n6960_t;wire n6961;wire n6961_t;wire n6962;wire n6962_t;wire n6963;wire n6963_t;wire n6964;wire n6964_t;wire n6965;wire n6965_t;wire n6966;wire n6966_t;wire n6967;wire n6967_t;wire n6968;wire n6968_t;wire n6969;wire n6969_t;wire n6970;wire n6970_t;wire n6971;wire n6971_t;wire n6972;wire n6972_t;wire n6973;wire n6973_t;wire n6974;wire n6974_t;wire n6975;wire n6975_t;wire n6976;wire n6976_t;wire n6977;wire n6977_t;wire n6978;wire n6978_t;wire n6979;wire n6979_t;wire n6980;wire n6980_t;wire n6981;wire n6981_t;wire n6982;wire n6982_t;wire n6983;wire n6983_t;wire n6984;wire n6984_t;wire n6985;wire n6985_t;wire n6986;wire n6986_t;wire n6987;wire n6987_t;wire n6988;wire n6988_t;wire n6989;wire n6989_t;wire n6990;wire n6990_t;wire n6991;wire n6991_t;wire n6992;wire n6992_t;wire n6993;wire n6993_t;wire n6994;wire n6994_t;wire n6995;wire n6995_t;wire n6996;wire n6996_t;wire n6997;wire n6997_t;wire n6998;wire n6998_t;wire n6999;wire n6999_t;wire n7000;wire n7000_t;wire n7001;wire n7001_t;wire n7002;wire n7002_t;wire n7003;wire n7003_t;wire n7004;wire n7004_t;wire n7005;wire n7005_t;wire n7006;wire n7006_t;wire n7007;wire n7007_t;wire n7008;wire n7008_t;wire n7009;wire n7009_t;wire n7010;wire n7010_t;wire n7011;wire n7011_t;wire n7012;wire n7012_t;wire n7013;wire n7013_t;wire n7014;wire n7014_t;wire n7015;wire n7015_t;wire n7016;wire n7016_t;wire n7017;wire n7017_t;wire n7018;wire n7018_t;wire n7019;wire n7019_t;wire n7020;wire n7020_t;wire n7021;wire n7021_t;wire n7022;wire n7022_t;wire n7023;wire n7023_t;wire n7024;wire n7024_t;wire n7025;wire n7025_t;wire n7026;wire n7026_t;wire n7027;wire n7027_t;wire n7028;wire n7028_t;wire n7029;wire n7029_t;wire n7030;wire n7030_t;wire n7031;wire n7031_t;wire n7032;wire n7032_t;wire n7033;wire n7033_t;wire n7034;wire n7034_t;wire n7035;wire n7035_t;wire n7036;wire n7036_t;wire n7037;wire n7037_t;wire n7038;wire n7038_t;wire n7039;wire n7039_t;wire n7040;wire n7040_t;wire n7041;wire n7041_t;wire n7042;wire n7042_t;wire n7043;wire n7043_t;wire n7044;wire n7044_t;wire n7045;wire n7045_t;wire n7046;wire n7046_t;wire n7047;wire n7047_t;wire n7048;wire n7048_t;wire n7049;wire n7049_t;wire n7050;wire n7050_t;wire n7051;wire n7051_t;wire n7052;wire n7052_t;wire n7053;wire n7053_t;wire n7054;wire n7054_t;wire n7055;wire n7055_t;wire n7056;wire n7056_t;wire n7057;wire n7057_t;wire n7058;wire n7058_t;wire n7059;wire n7059_t;wire n7060;wire n7060_t;wire n7061;wire n7061_t;wire n7062;wire n7062_t;wire n7063;wire n7063_t;wire n7064;wire n7064_t;wire n7065;wire n7065_t;wire n7066;wire n7066_t;wire n7067;wire n7067_t;wire n7068;wire n7068_t;wire n7069;wire n7069_t;wire n7070;wire n7070_t;wire n7071;wire n7071_t;wire n7072;wire n7072_t;wire n7073;wire n7073_t;wire n7074;wire n7074_t;wire n7075;wire n7075_t;wire n7076;wire n7076_t;wire n7077;wire n7077_t;wire n7078;wire n7078_t;wire n7079;wire n7079_t;wire n7080;wire n7080_t;wire n7081;wire n7081_t;wire n7082;wire n7082_t;wire n7083;wire n7083_t;wire n7084;wire n7084_t;wire n7085;wire n7085_t;wire n7086;wire n7086_t;wire n7087;wire n7087_t;wire n7088;wire n7088_t;wire n7089;wire n7089_t;wire n7090;wire n7090_t;wire n7091;wire n7091_t;wire n7092;wire n7092_t;wire n7093;wire n7093_t;wire n7094;wire n7094_t;wire n7095;wire n7095_t;wire n7096;wire n7096_t;wire n7097;wire n7097_t;wire n7098;wire n7098_t;wire n7099;wire n7099_t;wire n7100;wire n7100_t;wire n7101;wire n7101_t;wire n7102;wire n7102_t;wire n7103;wire n7103_t;wire n7104;wire n7104_t;wire n7105;wire n7105_t;wire n7106;wire n7106_t;wire n7107;wire n7107_t;wire n7108;wire n7108_t;wire n7109;wire n7109_t;wire n7110;wire n7110_t;wire n7111;wire n7111_t;wire n7112;wire n7112_t;wire n7113;wire n7113_t;wire n7114;wire n7114_t;wire n7115;wire n7115_t;wire n7116;wire n7116_t;wire n7117;wire n7117_t;wire n7118;wire n7118_t;wire n7119;wire n7119_t;wire n7120;wire n7120_t;wire n7121;wire n7121_t;wire n7122;wire n7122_t;wire n7123;wire n7123_t;wire n7124;wire n7124_t;wire n7125;wire n7125_t;wire n7126;wire n7126_t;wire n7127;wire n7127_t;wire n7128;wire n7128_t;wire n7129;wire n7129_t;wire n7130;wire n7130_t;wire n7131;wire n7131_t;wire n7132;wire n7132_t;wire n7133;wire n7133_t;wire n7134;wire n7134_t;wire n7135;wire n7135_t;wire n7136;wire n7136_t;wire n7137;wire n7137_t;wire n7138;wire n7138_t;wire n7139;wire n7139_t;wire n7140;wire n7140_t;wire n7141;wire n7141_t;wire n7142;wire n7142_t;wire n7143;wire n7143_t;wire n7144;wire n7144_t;wire n7145;wire n7145_t;wire n7146;wire n7146_t;wire n7147;wire n7147_t;wire n7148;wire n7148_t;wire n7149;wire n7149_t;wire n7150;wire n7150_t;wire n7151;wire n7151_t;wire n7152;wire n7152_t;wire n7153;wire n7153_t;wire n7154;wire n7154_t;wire n7155;wire n7155_t;wire n7156;wire n7156_t;wire n7157;wire n7157_t;wire n7158;wire n7158_t;wire n7159;wire n7159_t;wire n7160;wire n7160_t;wire n7161;wire n7161_t;wire n7162;wire n7162_t;wire n7163;wire n7163_t;wire n7164;wire n7164_t;wire n7165;wire n7165_t;wire n7166;wire n7166_t;wire n7167;wire n7167_t;wire n7168;wire n7168_t;wire n7169;wire n7169_t;wire n7170;wire n7170_t;wire n7171;wire n7171_t;wire n7172;wire n7172_t;wire n7173;wire n7173_t;wire n7174;wire n7174_t;wire n7175;wire n7175_t;wire n7176;wire n7176_t;wire n7177;wire n7177_t;wire n7178;wire n7178_t;wire n7179;wire n7179_t;wire n7180;wire n7180_t;wire n7181;wire n7181_t;wire n7182;wire n7182_t;wire n7183;wire n7183_t;wire n7184;wire n7184_t;wire n7185;wire n7185_t;wire n7186;wire n7186_t;wire n7187;wire n7187_t;wire n7188;wire n7188_t;wire n7189;wire n7189_t;wire n7190;wire n7190_t;wire n7191;wire n7191_t;wire n7192;wire n7192_t;wire n7193;wire n7193_t;wire n7194;wire n7194_t;wire n7195;wire n7195_t;wire n7196;wire n7196_t;wire n7197;wire n7197_t;wire n7198;wire n7198_t;wire n7199;wire n7199_t;wire n7200;wire n7200_t;wire n7201;wire n7201_t;wire n7202;wire n7202_t;wire n7203;wire n7203_t;wire n7204;wire n7204_t;wire n7205;wire n7205_t;wire n7206;wire n7206_t;wire n7207;wire n7207_t;wire n7208;wire n7208_t;wire n7209;wire n7209_t;wire n7210;wire n7210_t;wire n7211;wire n7211_t;wire n7212;wire n7212_t;wire n7213;wire n7213_t;wire n7214;wire n7214_t;wire n7215;wire n7215_t;wire n7216;wire n7216_t;wire n7217;wire n7217_t;wire n7218;wire n7218_t;wire n7219;wire n7219_t;wire n7220;wire n7220_t;wire n7221;wire n7221_t;wire n7222;wire n7222_t;wire n7223;wire n7223_t;wire n7224;wire n7224_t;wire n7225;wire n7225_t;wire n7226;wire n7226_t;wire n7227;wire n7227_t;wire n7228;wire n7228_t;wire n7229;wire n7229_t;wire n7230;wire n7230_t;wire n7231;wire n7231_t;wire n7232;wire n7232_t;wire n7233;wire n7233_t;wire n7234;wire n7234_t;wire n7235;wire n7235_t;wire n7236;wire n7236_t;wire n7237;wire n7237_t;wire n7238;wire n7238_t;wire n7239;wire n7239_t;wire n7240;wire n7240_t;wire n7241;wire n7241_t;wire n7242;wire n7242_t;wire n7243;wire n7243_t;wire n7244;wire n7244_t;wire n7245;wire n7245_t;wire n7246;wire n7246_t;wire n7247;wire n7247_t;wire n7248;wire n7248_t;wire n7249;wire n7249_t;wire n7250;wire n7250_t;wire n7251;wire n7251_t;wire n7252;wire n7252_t;wire n7253;wire n7253_t;wire n7254;wire n7254_t;wire n7255;wire n7255_t;wire n7256;wire n7256_t;wire n7257;wire n7257_t;wire n7258;wire n7258_t;wire n7259;wire n7259_t;wire n7260;wire n7260_t;wire n7261;wire n7261_t;wire n7262;wire n7262_t;wire n7263;wire n7263_t;wire n7264;wire n7264_t;wire n7265;wire n7265_t;wire n7266;wire n7266_t;wire n7267;wire n7267_t;wire n7268;wire n7268_t;wire n7269;wire n7269_t;wire n7270;wire n7270_t;wire n7271;wire n7271_t;wire n7272;wire n7272_t;wire n7273;wire n7273_t;wire n7274;wire n7274_t;wire n7275;wire n7275_t;wire n7276;wire n7276_t;wire n7277;wire n7277_t;wire n7278;wire n7278_t;wire n7279;wire n7279_t;wire n7280;wire n7280_t;wire n7281;wire n7281_t;wire n7282;wire n7282_t;wire n7283;wire n7283_t;wire n7284;wire n7284_t;wire n7285;wire n7285_t;wire n7286;wire n7286_t;wire n7287;wire n7287_t;wire n7288;wire n7288_t;wire n7289;wire n7289_t;wire n7290;wire n7290_t;wire n7291;wire n7291_t;wire n7292;wire n7292_t;wire n7293;wire n7293_t;wire n7294;wire n7294_t;wire n7295;wire n7295_t;wire n7296;wire n7296_t;wire n7297;wire n7297_t;wire n7298;wire n7298_t;wire n7299;wire n7299_t;wire n7300;wire n7300_t;wire n7301;wire n7301_t;wire n7302;wire n7302_t;wire n7303;wire n7303_t;wire n7304;wire n7304_t;wire n7305;wire n7305_t;wire n7306;wire n7306_t;wire n7307;wire n7307_t;wire n7308;wire n7308_t;wire n7309;wire n7309_t;wire n7310;wire n7310_t;wire n7311;wire n7311_t;wire n7312;wire n7312_t;wire n7313;wire n7313_t;wire n7314;wire n7314_t;wire n7315;wire n7315_t;wire n7316;wire n7316_t;wire n7317;wire n7317_t;wire n7318;wire n7318_t;wire n7319;wire n7319_t;wire n7320;wire n7320_t;wire n7321;wire n7321_t;wire n7322;wire n7322_t;wire n7323;wire n7323_t;wire n7324;wire n7324_t;wire n7325;wire n7325_t;wire n7326;wire n7326_t;wire n7327;wire n7327_t;wire n7328;wire n7328_t;wire n7329;wire n7329_t;wire n7330;wire n7330_t;wire n7331;wire n7331_t;wire n7332;wire n7332_t;wire n7333;wire n7333_t;wire n7334;wire n7334_t;wire n7335;wire n7335_t;wire n7336;wire n7336_t;wire n7337;wire n7337_t;wire n7338;wire n7338_t;wire n7339;wire n7339_t;wire n7340;wire n7340_t;wire n7341;wire n7341_t;wire n7342;wire n7342_t;wire n7343;wire n7343_t;wire n7344;wire n7344_t;wire n7345;wire n7345_t;wire n7346;wire n7346_t;wire n7347;wire n7347_t;wire n7348;wire n7348_t;wire n7349;wire n7349_t;wire n7350;wire n7350_t;wire n7351;wire n7351_t;wire n7352;wire n7352_t;wire n7353;wire n7353_t;wire n7354;wire n7354_t;wire n7355;wire n7355_t;wire n7356;wire n7356_t;wire n7357;wire n7357_t;wire n7358;wire n7358_t;wire n7359;wire n7359_t;wire n7360;wire n7360_t;wire n7361;wire n7361_t;wire n7362;wire n7362_t;wire n7363;wire n7363_t;wire n7364;wire n7364_t;wire n7365;wire n7365_t;wire n7366;wire n7366_t;wire n7367;wire n7367_t;wire n7368;wire n7368_t;wire n7369;wire n7369_t;wire n7370;wire n7370_t;wire n7371;wire n7371_t;wire n7372;wire n7372_t;wire n7373;wire n7373_t;wire n7374;wire n7374_t;wire n7375;wire n7375_t;wire n7376;wire n7376_t;wire n7377;wire n7377_t;wire n7378;wire n7378_t;wire n7379;wire n7379_t;wire n7380;wire n7380_t;wire n7381;wire n7381_t;wire n7382;wire n7382_t;wire n7383;wire n7383_t;wire n7384;wire n7384_t;wire n7385;wire n7385_t;wire n7386;wire n7386_t;wire n7387;wire n7387_t;wire n7388;wire n7388_t;wire n7389;wire n7389_t;wire n7390;wire n7390_t;wire n7391;wire n7391_t;wire n7392;wire n7392_t;wire n7393;wire n7393_t;wire n7394;wire n7394_t;wire n7395;wire n7395_t;wire n7396;wire n7396_t;wire n7397;wire n7397_t;wire n7398;wire n7398_t;wire n7399;wire n7399_t;wire n7400;wire n7400_t;wire n7401;wire n7401_t;wire n7402;wire n7402_t;wire n7403;wire n7403_t;wire n7404;wire n7404_t;wire n7405;wire n7405_t;wire n7406;wire n7406_t;wire n7407;wire n7407_t;wire n7408;wire n7408_t;wire n7409;wire n7409_t;wire n7410;wire n7410_t;wire n7411;wire n7411_t;wire n7412;wire n7412_t;wire n7413;wire n7413_t;wire n7414;wire n7414_t;wire n7415;wire n7415_t;wire n7416;wire n7416_t;wire n7417;wire n7417_t;wire n7418;wire n7418_t;wire n7419;wire n7419_t;wire n7420;wire n7420_t;wire n7421;wire n7421_t;wire n7422;wire n7422_t;wire n7423;wire n7423_t;wire n7424;wire n7424_t;wire n7425;wire n7425_t;wire n7426;wire n7426_t;wire n7427;wire n7427_t;wire n7428;wire n7428_t;wire n7429;wire n7429_t;wire n7430;wire n7430_t;wire n7431;wire n7431_t;wire n7432;wire n7432_t;wire n7433;wire n7433_t;wire n7434;wire n7434_t;wire n7435;wire n7435_t;wire n7436;wire n7436_t;wire n7437;wire n7437_t;wire n7438;wire n7438_t;wire n7439;wire n7439_t;wire n7440;wire n7440_t;wire n7441;wire n7441_t;wire n7442;wire n7442_t;wire n7443;wire n7443_t;wire n7444;wire n7444_t;wire n7445;wire n7445_t;wire n7446;wire n7446_t;wire n7447;wire n7447_t;wire n7448;wire n7448_t;wire n7449;wire n7449_t;wire n7450;wire n7450_t;wire n7451;wire n7451_t;wire n7452;wire n7452_t;wire n7453;wire n7453_t;wire n7454;wire n7454_t;wire n7455;wire n7455_t;wire n7456;wire n7456_t;wire n7457;wire n7457_t;wire n7458;wire n7458_t;wire n7459;wire n7459_t;wire n7460;wire n7460_t;wire n7461;wire n7461_t;wire n7462;wire n7462_t;wire n7463;wire n7463_t;wire n7464;wire n7464_t;wire n7465;wire n7465_t;wire n7466;wire n7466_t;wire n7467;wire n7467_t;wire n7468;wire n7468_t;wire n7469;wire n7469_t;wire n7470;wire n7470_t;wire n7471;wire n7471_t;wire n7472;wire n7472_t;wire n7473;wire n7473_t;wire n7474;wire n7474_t;wire n7475;wire n7475_t;wire n7476;wire n7476_t;wire n7477;wire n7477_t;wire n7478;wire n7478_t;wire n7479;wire n7479_t;wire n7480;wire n7480_t;wire n7481;wire n7481_t;wire n7482;wire n7482_t;wire n7483;wire n7483_t;wire n7484;wire n7484_t;wire n7485;wire n7485_t;wire n7486;wire n7486_t;wire n7487;wire n7487_t;wire n7488;wire n7488_t;wire n7489;wire n7489_t;wire n7490;wire n7490_t;wire n7491;wire n7491_t;wire n7492;wire n7492_t;wire n7493;wire n7493_t;wire n7494;wire n7494_t;wire n7495;wire n7495_t;wire n7496;wire n7496_t;wire n7497;wire n7497_t;wire n7498;wire n7498_t;wire n7499;wire n7499_t;wire n7500;wire n7500_t;wire n7501;wire n7501_t;wire n7502;wire n7502_t;wire n7503;wire n7503_t;wire n7504;wire n7504_t;wire n7505;wire n7505_t;wire n7506;wire n7506_t;wire n7507;wire n7507_t;wire n7508;wire n7508_t;wire n7509;wire n7509_t;wire n7510;wire n7510_t;wire n7511;wire n7511_t;wire n7512;wire n7512_t;wire n7513;wire n7513_t;wire n7514;wire n7514_t;wire n7515;wire n7515_t;wire n7516;wire n7516_t;wire n7517;wire n7517_t;wire n7518;wire n7518_t;wire n7519;wire n7519_t;wire n7520;wire n7520_t;wire n7521;wire n7521_t;wire n7522;wire n7522_t;wire n7523;wire n7523_t;wire n7524;wire n7524_t;wire n7525;wire n7525_t;wire n7526;wire n7526_t;wire n7527;wire n7527_t;wire n7528;wire n7528_t;wire n7529;wire n7529_t;wire n7530;wire n7530_t;wire n7531;wire n7531_t;wire n7532;wire n7532_t;wire n7533;wire n7533_t;wire n7534;wire n7534_t;wire n7535;wire n7535_t;wire n7536;wire n7536_t;wire n7537;wire n7537_t;wire n7538;wire n7538_t;wire n7539;wire n7539_t;wire n7540;wire n7540_t;wire n7541;wire n7541_t;wire n7542;wire n7542_t;wire n7543;wire n7543_t;wire n7544;wire n7544_t;wire n7545;wire n7545_t;wire n7546;wire n7546_t;wire n7547;wire n7547_t;wire n7548;wire n7548_t;wire n7549;wire n7549_t;wire n7550;wire n7550_t;wire n7551;wire n7551_t;wire n7552;wire n7552_t;wire n7553;wire n7553_t;wire n7554;wire n7554_t;wire n7555;wire n7555_t;wire n7556;wire n7556_t;wire n7557;wire n7557_t;wire n7558;wire n7558_t;wire n7559;wire n7559_t;wire n7560;wire n7560_t;wire n7561;wire n7561_t;wire n7562;wire n7562_t;wire n7563;wire n7563_t;wire n7564;wire n7564_t;wire n7565;wire n7565_t;wire n7566;wire n7566_t;wire n7567;wire n7567_t;wire n7568;wire n7568_t;wire n7569;wire n7569_t;wire n7570;wire n7570_t;wire n7571;wire n7571_t;wire n7572;wire n7572_t;wire n7573;wire n7573_t;wire n7574;wire n7574_t;wire n7575;wire n7575_t;wire n7576;wire n7576_t;wire n7577;wire n7577_t;wire n7578;wire n7578_t;wire n7579;wire n7579_t;wire n7580;wire n7580_t;wire n7581;wire n7581_t;wire n7582;wire n7582_t;wire n7583;wire n7583_t;wire n7584;wire n7584_t;wire n7585;wire n7585_t;wire n7586;wire n7586_t;wire n7587;wire n7587_t;wire n7588;wire n7588_t;wire n7589;wire n7589_t;wire n7590;wire n7590_t;wire n7591;wire n7591_t;wire n7592;wire n7592_t;wire n7593;wire n7593_t;wire n7594;wire n7594_t;wire n7595;wire n7595_t;wire n7596;wire n7596_t;wire n7597;wire n7597_t;wire n7598;wire n7598_t;wire n7599;wire n7599_t;wire n7600;wire n7600_t;wire n7601;wire n7601_t;wire n7602;wire n7602_t;wire n7603;wire n7603_t;wire n7604;wire n7604_t;wire n7605;wire n7605_t;wire n7606;wire n7606_t;wire n7607;wire n7607_t;wire n7608;wire n7608_t;wire n7609;wire n7609_t;wire n7610;wire n7610_t;wire n7611;wire n7611_t;wire n7612;wire n7612_t;wire n7613;wire n7613_t;wire n7614;wire n7614_t;wire n7615;wire n7615_t;wire n7616;wire n7616_t;wire n7617;wire n7617_t;wire n7618;wire n7618_t;wire n7619;wire n7619_t;wire n7620;wire n7620_t;wire n7621;wire n7621_t;wire n7622;wire n7622_t;wire n7623;wire n7623_t;wire n7624;wire n7624_t;wire n7625;wire n7625_t;wire n7626;wire n7626_t;wire n7627;wire n7627_t;wire n7628;wire n7628_t;wire n7629;wire n7629_t;wire n7630;wire n7630_t;wire n7631;wire n7631_t;wire n7632;wire n7632_t;wire n7633;wire n7633_t;wire n7634;wire n7634_t;wire n7635;wire n7635_t;wire n7636;wire n7636_t;wire n7637;wire n7637_t;wire n7638;wire n7638_t;wire n7639;wire n7639_t;wire n7640;wire n7640_t;wire n7641;wire n7641_t;wire n7642;wire n7642_t;wire n7643;wire n7643_t;wire n7644;wire n7644_t;wire n7645;wire n7645_t;wire n7646;wire n7646_t;wire n7647;wire n7647_t;wire n7648;wire n7648_t;wire n7649;wire n7649_t;wire n7650;wire n7650_t;wire n7651;wire n7651_t;wire n7652;wire n7652_t;wire n7653;wire n7653_t;wire n7654;wire n7654_t;wire n7655;wire n7655_t;wire n7656;wire n7656_t;wire n7657;wire n7657_t;wire n7658;wire n7658_t;wire n7659;wire n7659_t;wire n7660;wire n7660_t;wire n7661;wire n7661_t;wire n7662;wire n7662_t;wire n7663;wire n7663_t;wire n7664;wire n7664_t;wire n7665;wire n7665_t;wire n7666;wire n7666_t;wire n7667;wire n7667_t;wire n7668;wire n7668_t;wire n7669;wire n7669_t;wire n7670;wire n7670_t;wire n7671;wire n7671_t;wire n7672;wire n7672_t;wire n7673;wire n7673_t;wire n7674;wire n7674_t;wire n7675;wire n7675_t;wire n7676;wire n7676_t;wire n7677;wire n7677_t;wire n7678;wire n7678_t;wire n7679;wire n7679_t;wire n7680;wire n7680_t;wire n7681;wire n7681_t;wire n7682;wire n7682_t;wire n7683;wire n7683_t;wire n7684;wire n7684_t;wire n7685;wire n7685_t;wire n7686;wire n7686_t;wire n7687;wire n7687_t;wire n7688;wire n7688_t;wire n7689;wire n7689_t;wire n7690;wire n7690_t;wire n7691;wire n7691_t;wire n7692;wire n7692_t;wire n7693;wire n7693_t;wire n7694;wire n7694_t;wire n7695;wire n7695_t;wire n7696;wire n7696_t;wire n7697;wire n7697_t;wire n7698;wire n7698_t;wire n7699;wire n7699_t;wire n7700;wire n7700_t;wire n7701;wire n7701_t;wire n7702;wire n7702_t;wire n7703;wire n7703_t;wire n7704;wire n7704_t;wire n7705;wire n7705_t;wire n7706;wire n7706_t;wire n7707;wire n7707_t;wire n7708;wire n7708_t;wire n7709;wire n7709_t;wire n7710;wire n7710_t;wire n7711;wire n7711_t;wire n7712;wire n7712_t;wire n7713;wire n7713_t;wire n7714;wire n7714_t;wire n7715;wire n7715_t;wire n7716;wire n7716_t;wire n7717;wire n7717_t;wire n7718;wire n7718_t;wire n7719;wire n7719_t;wire n7720;wire n7720_t;wire n7721;wire n7721_t;wire n7722;wire n7722_t;wire n7723;wire n7723_t;wire n7724;wire n7724_t;wire n7725;wire n7725_t;wire n7726;wire n7726_t;wire n7727;wire n7727_t;wire n7728;wire n7728_t;wire n7729;wire n7729_t;wire n7730;wire n7730_t;wire n7731;wire n7731_t;wire n7732;wire n7732_t;wire n7733;wire n7733_t;wire n7734;wire n7734_t;wire n7735;wire n7735_t;wire n7736;wire n7736_t;wire n7737;wire n7737_t;wire n7738;wire n7738_t;wire n7739;wire n7739_t;wire n7740;wire n7740_t;wire n7741;wire n7741_t;wire n7742;wire n7742_t;wire n7743;wire n7743_t;wire n7744;wire n7744_t;wire n7745;wire n7745_t;wire n7746;wire n7746_t;wire n7747;wire n7747_t;wire n7748;wire n7748_t;wire n7749;wire n7749_t;wire n7750;wire n7750_t;wire n7751;wire n7751_t;wire n7752;wire n7752_t;wire n7753;wire n7753_t;wire n7754;wire n7754_t;wire n7755;wire n7755_t;wire n7756;wire n7756_t;wire n7757;wire n7757_t;wire n7758;wire n7758_t;wire n7759;wire n7759_t;wire n7760;wire n7760_t;wire n7761;wire n7761_t;wire n7762;wire n7762_t;wire n7763;wire n7763_t;wire n7764;wire n7764_t;wire n7765;wire n7765_t;wire n7766;wire n7766_t;wire n7767;wire n7767_t;wire n7768;wire n7768_t;wire n7769;wire n7769_t;wire n7770;wire n7770_t;wire n7771;wire n7771_t;wire n7772;wire n7772_t;wire n7773;wire n7773_t;wire n7774;wire n7774_t;wire n7775;wire n7775_t;wire n7776;wire n7776_t;wire n7777;wire n7777_t;wire n7778;wire n7778_t;wire n7779;wire n7779_t;wire n7780;wire n7780_t;wire n7781;wire n7781_t;wire n7782;wire n7782_t;wire n7783;wire n7783_t;wire n7784;wire n7784_t;wire n7785;wire n7785_t;wire n7786;wire n7786_t;wire n7787;wire n7787_t;wire n7788;wire n7788_t;wire n7789;wire n7789_t;wire n7790;wire n7790_t;wire n7791;wire n7791_t;wire n7792;wire n7792_t;wire n7793;wire n7793_t;wire n7794;wire n7794_t;wire n7795;wire n7795_t;wire n7796;wire n7796_t;wire n7797;wire n7797_t;wire n7798;wire n7798_t;wire n7799;wire n7799_t;wire n7800;wire n7800_t;wire n7801;wire n7801_t;wire n7802;wire n7802_t;wire n7803;wire n7803_t;wire n7804;wire n7804_t;wire n7805;wire n7805_t;wire n7806;wire n7806_t;wire n7807;wire n7807_t;wire n7808;wire n7808_t;wire n7809;wire n7809_t;wire n7810;wire n7810_t;wire n7811;wire n7811_t;wire n7812;wire n7812_t;wire n7813;wire n7813_t;wire n7814;wire n7814_t;wire n7815;wire n7815_t;wire n7816;wire n7816_t;wire n7817;wire n7817_t;wire n7818;wire n7818_t;wire n7819;wire n7819_t;wire n7820;wire n7820_t;wire n7821;wire n7821_t;wire n7822;wire n7822_t;wire n7823;wire n7823_t;wire n7824;wire n7824_t;wire n7825;wire n7825_t;wire n7826;wire n7826_t;wire n7827;wire n7827_t;wire n7828;wire n7828_t;wire n7829;wire n7829_t;wire n7830;wire n7830_t;wire n7831;wire n7831_t;wire n7832;wire n7832_t;wire n7833;wire n7833_t;wire n7834;wire n7834_t;wire n7835;wire n7835_t;wire n7836;wire n7836_t;wire n7837;wire n7837_t;wire n7838;wire n7838_t;wire n7839;wire n7839_t;wire n7840;wire n7840_t;wire n7841;wire n7841_t;wire n7842;wire n7842_t;wire n7843;wire n7843_t;wire n7844;wire n7844_t;wire n7845;wire n7845_t;wire n7846;wire n7846_t;wire n7847;wire n7847_t;wire n7848;wire n7848_t;wire n7849;wire n7849_t;wire n7850;wire n7850_t;wire n7851;wire n7851_t;wire n7852;wire n7852_t;wire n7853;wire n7853_t;wire n7854;wire n7854_t;wire n7855;wire n7855_t;wire n7856;wire n7856_t;wire n7857;wire n7857_t;wire n7858;wire n7858_t;wire n7859;wire n7859_t;wire n7860;wire n7860_t;wire n7861;wire n7861_t;wire n7862;wire n7862_t;wire n7863;wire n7863_t;wire n7864;wire n7864_t;wire n7865;wire n7865_t;wire n7866;wire n7866_t;wire n7867;wire n7867_t;wire n7868;wire n7868_t;wire n7869;wire n7869_t;wire n7870;wire n7870_t;wire n7871;wire n7871_t;wire n7872;wire n7872_t;wire n7873;wire n7873_t;wire n7874;wire n7874_t;wire n7875;wire n7875_t;wire n7876;wire n7876_t;wire n7877;wire n7877_t;wire n7878;wire n7878_t;wire n7879;wire n7879_t;wire n7880;wire n7880_t;wire n7881;wire n7881_t;wire n7882;wire n7882_t;wire n7883;wire n7883_t;wire n7884;wire n7884_t;wire n7885;wire n7885_t;wire n7886;wire n7886_t;wire n7887;wire n7887_t;wire n7888;wire n7888_t;wire n7889;wire n7889_t;wire n7890;wire n7890_t;wire n7891;wire n7891_t;wire n7892;wire n7892_t;wire n7893;wire n7893_t;wire n7894;wire n7894_t;wire n7895;wire n7895_t;wire n7896;wire n7896_t;wire n7897;wire n7897_t;wire n7898;wire n7898_t;wire n7899;wire n7899_t;wire n7900;wire n7900_t;wire n7901;wire n7901_t;wire n7902;wire n7902_t;wire n7903;wire n7903_t;wire n7904;wire n7904_t;wire n7905;wire n7905_t;wire n7906;wire n7906_t;wire n7907;wire n7907_t;wire n7908;wire n7908_t;wire n7909;wire n7909_t;wire n7910;wire n7910_t;wire n7911;wire n7911_t;wire n7912;wire n7912_t;wire n7913;wire n7913_t;wire n7914;wire n7914_t;wire n7915;wire n7915_t;wire n7916;wire n7916_t;wire n7917;wire n7917_t;wire n7918;wire n7918_t;wire n7919;wire n7919_t;wire n7920;wire n7920_t;wire n7921;wire n7921_t;wire n7922;wire n7922_t;wire n7923;wire n7923_t;wire n7924;wire n7924_t;wire n7925;wire n7925_t;wire n7926;wire n7926_t;wire n7927;wire n7927_t;wire n7928;wire n7928_t;wire n7929;wire n7929_t;wire n7930;wire n7930_t;wire n7931;wire n7931_t;wire n7932;wire n7932_t;wire n7933;wire n7933_t;wire n7934;wire n7934_t;wire n7935;wire n7935_t;wire n7936;wire n7936_t;wire n7937;wire n7937_t;wire n7938;wire n7938_t;wire n7939;wire n7939_t;wire n7940;wire n7940_t;wire n7941;wire n7941_t;wire n7942;wire n7942_t;wire n7943;wire n7943_t;wire n7944;wire n7944_t;wire n7945;wire n7945_t;wire n7946;wire n7946_t;wire n7947;wire n7947_t;wire n7948;wire n7948_t;wire n7949;wire n7949_t;wire n7950;wire n7950_t;wire n7951;wire n7951_t;wire n7952;wire n7952_t;wire n7953;wire n7953_t;wire n7954;wire n7954_t;wire n7955;wire n7955_t;wire n7956;wire n7956_t;wire n7957;wire n7957_t;wire n7958;wire n7958_t;wire n7959;wire n7959_t;wire n7960;wire n7960_t;wire n7961;wire n7961_t;wire n7962;wire n7962_t;wire n7963;wire n7963_t;wire n7964;wire n7964_t;wire n7965;wire n7965_t;wire n7966;wire n7966_t;wire n7967;wire n7967_t;wire n7968;wire n7968_t;wire n7969;wire n7969_t;wire n7970;wire n7970_t;wire n7971;wire n7971_t;wire n7972;wire n7972_t;wire n7973;wire n7973_t;wire n7974;wire n7974_t;wire n7975;wire n7975_t;wire n7976;wire n7976_t;wire n7977;wire n7977_t;wire n7978;wire n7978_t;wire n7979;wire n7979_t;wire n7980;wire n7980_t;wire n7981;wire n7981_t;wire n7982;wire n7982_t;wire n7983;wire n7983_t;wire n7984;wire n7984_t;wire n7985;wire n7985_t;wire n7986;wire n7986_t;wire n7987;wire n7987_t;wire n7988;wire n7988_t;wire n7989;wire n7989_t;wire n7990;wire n7990_t;wire n7991;wire n7991_t;wire n7992;wire n7992_t;wire n7993;wire n7993_t;wire n7994;wire n7994_t;
  wire Trigger_en10_0;wire Trigger_en10_0_t;wire troj10_0n1;wire troj10_0n1_t;wire troj10_0n2;wire troj10_0n2_t;wire troj10_0n3;wire troj10_0n3_t;wire troj10_0n4;wire troj10_0n4_t;wire troj10_0n5;wire troj10_0n5_t;wire troj10_0n6;wire troj10_0n6_t;wire tempn3869;wire tempn3869_t;wire Trigger_en10_1;wire Trigger_en10_1_t;wire troj10_1n1;wire troj10_1n1_t;wire troj10_1n2;wire troj10_1n2_t;wire troj10_1n3;wire troj10_1n3_t;wire troj10_1n4;wire troj10_1n4_t;wire tempn2493;wire tempn2493_t;
  assign test_so = CRC_OUT_1_31;
  assign test_so_t = CRC_OUT_1_31_t;

  nor2s3
  U1
  (
    .DIN1(n4997),
    .DIN1_t(n4997_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX9949),
    .Q_t(WX9949_t)
  );


  nor2s3
  U2
  (
    .DIN1(n5001),
    .DIN1_t(n5001_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX9947),
    .Q_t(WX9947_t)
  );


  nor2s3
  U3
  (
    .DIN1(n5005),
    .DIN1_t(n5005_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX9945),
    .Q_t(WX9945_t)
  );


  nor2s3
  U4
  (
    .DIN1(n5009),
    .DIN1_t(n5009_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX9943),
    .Q_t(WX9943_t)
  );


  nor2s3
  U5
  (
    .DIN1(n5013),
    .DIN1_t(n5013_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX9941),
    .Q_t(WX9941_t)
  );


  nor2s3
  U6
  (
    .DIN1(n5017),
    .DIN1_t(n5017_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9939),
    .Q_t(WX9939_t)
  );


  nor2s3
  U7
  (
    .DIN1(n5021),
    .DIN1_t(n5021_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9937),
    .Q_t(WX9937_t)
  );


  nor2s3
  U8
  (
    .DIN1(n5025),
    .DIN1_t(n5025_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9935),
    .Q_t(WX9935_t)
  );


  nor2s3
  U9
  (
    .DIN1(n5029),
    .DIN1_t(n5029_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9933),
    .Q_t(WX9933_t)
  );


  nor2s3
  U10
  (
    .DIN1(n5033),
    .DIN1_t(n5033_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9931),
    .Q_t(WX9931_t)
  );


  nor2s3
  U11
  (
    .DIN1(n5037),
    .DIN1_t(n5037_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9929),
    .Q_t(WX9929_t)
  );


  nor2s3
  U12
  (
    .DIN1(n5041),
    .DIN1_t(n5041_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9927),
    .Q_t(WX9927_t)
  );


  nor2s3
  U13
  (
    .DIN1(n5045),
    .DIN1_t(n5045_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9925),
    .Q_t(WX9925_t)
  );


  nor2s3
  U14
  (
    .DIN1(n5049),
    .DIN1_t(n5049_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9923),
    .Q_t(WX9923_t)
  );


  nor2s3
  U15
  (
    .DIN1(n5053),
    .DIN1_t(n5053_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9921),
    .Q_t(WX9921_t)
  );


  nor2s3
  U16
  (
    .DIN1(n5057),
    .DIN1_t(n5057_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9919),
    .Q_t(WX9919_t)
  );


  nor2s3
  U17
  (
    .DIN1(n5061),
    .DIN1_t(n5061_t),
    .DIN2(n6744),
    .DIN2_t(n6744_t),
    .Q(WX9917),
    .Q_t(WX9917_t)
  );


  nor2s3
  U18
  (
    .DIN1(n5065),
    .DIN1_t(n5065_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9915),
    .Q_t(WX9915_t)
  );


  nor2s3
  U19
  (
    .DIN1(n5069),
    .DIN1_t(n5069_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9913),
    .Q_t(WX9913_t)
  );


  nor2s3
  U20
  (
    .DIN1(n5073),
    .DIN1_t(n5073_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9911),
    .Q_t(WX9911_t)
  );


  nor2s3
  U21
  (
    .DIN1(n5077),
    .DIN1_t(n5077_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9909),
    .Q_t(WX9909_t)
  );


  nor2s3
  U22
  (
    .DIN1(n5081),
    .DIN1_t(n5081_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9907),
    .Q_t(WX9907_t)
  );


  nor2s3
  U23
  (
    .DIN1(n5085),
    .DIN1_t(n5085_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9905),
    .Q_t(WX9905_t)
  );


  nor2s3
  U24
  (
    .DIN1(n5089),
    .DIN1_t(n5089_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9903),
    .Q_t(WX9903_t)
  );


  nor2s3
  U25
  (
    .DIN1(n5093),
    .DIN1_t(n5093_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9901),
    .Q_t(WX9901_t)
  );


  nor2s3
  U26
  (
    .DIN1(n5097),
    .DIN1_t(n5097_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9899),
    .Q_t(WX9899_t)
  );


  nor2s3
  U27
  (
    .DIN1(n5101),
    .DIN1_t(n5101_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9897),
    .Q_t(WX9897_t)
  );


  nor2s3
  U28
  (
    .DIN1(n5105),
    .DIN1_t(n5105_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9895),
    .Q_t(WX9895_t)
  );


  nor2s3
  U29
  (
    .DIN1(n5109),
    .DIN1_t(n5109_t),
    .DIN2(n6743),
    .DIN2_t(n6743_t),
    .Q(WX9893),
    .Q_t(WX9893_t)
  );


  nor2s3
  U30
  (
    .DIN1(n5113),
    .DIN1_t(n5113_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9891),
    .Q_t(WX9891_t)
  );


  nor2s3
  U31
  (
    .DIN1(n5117),
    .DIN1_t(n5117_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9889),
    .Q_t(WX9889_t)
  );


  nor2s3
  U32
  (
    .DIN1(n5121),
    .DIN1_t(n5121_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9887),
    .Q_t(WX9887_t)
  );


  nor2s3
  U33
  (
    .DIN1(n4996),
    .DIN1_t(n4996_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9885),
    .Q_t(WX9885_t)
  );


  nor2s3
  U34
  (
    .DIN1(n5000),
    .DIN1_t(n5000_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9883),
    .Q_t(WX9883_t)
  );


  nor2s3
  U35
  (
    .DIN1(n5004),
    .DIN1_t(n5004_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9881),
    .Q_t(WX9881_t)
  );


  nor2s3
  U36
  (
    .DIN1(n5008),
    .DIN1_t(n5008_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9879),
    .Q_t(WX9879_t)
  );


  nor2s3
  U37
  (
    .DIN1(n5012),
    .DIN1_t(n5012_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9877),
    .Q_t(WX9877_t)
  );


  nor2s3
  U38
  (
    .DIN1(n5016),
    .DIN1_t(n5016_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9875),
    .Q_t(WX9875_t)
  );


  nor2s3
  U39
  (
    .DIN1(n5020),
    .DIN1_t(n5020_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9873),
    .Q_t(WX9873_t)
  );


  nor2s3
  U40
  (
    .DIN1(n5024),
    .DIN1_t(n5024_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9871),
    .Q_t(WX9871_t)
  );


  nor2s3
  U41
  (
    .DIN1(n5028),
    .DIN1_t(n5028_t),
    .DIN2(n6742),
    .DIN2_t(n6742_t),
    .Q(WX9869),
    .Q_t(WX9869_t)
  );


  nor2s3
  U42
  (
    .DIN1(n5032),
    .DIN1_t(n5032_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9867),
    .Q_t(WX9867_t)
  );


  nor2s3
  U43
  (
    .DIN1(n5036),
    .DIN1_t(n5036_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9865),
    .Q_t(WX9865_t)
  );


  nor2s3
  U44
  (
    .DIN1(n5040),
    .DIN1_t(n5040_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9863),
    .Q_t(WX9863_t)
  );


  nor2s3
  U45
  (
    .DIN1(n5044),
    .DIN1_t(n5044_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9861),
    .Q_t(WX9861_t)
  );


  nor2s3
  U46
  (
    .DIN1(n5048),
    .DIN1_t(n5048_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9859),
    .Q_t(WX9859_t)
  );


  nor2s3
  U47
  (
    .DIN1(n5052),
    .DIN1_t(n5052_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9857),
    .Q_t(WX9857_t)
  );


  nor2s3
  U48
  (
    .DIN1(n5056),
    .DIN1_t(n5056_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9855),
    .Q_t(WX9855_t)
  );


  and2s3
  U49
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5060),
    .DIN2_t(n5060_t),
    .Q(WX9853),
    .Q_t(WX9853_t)
  );


  and2s3
  U50
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5064),
    .DIN2_t(n5064_t),
    .Q(WX9851),
    .Q_t(WX9851_t)
  );


  and2s3
  U51
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5068),
    .DIN2_t(n5068_t),
    .Q(WX9849),
    .Q_t(WX9849_t)
  );


  and2s3
  U52
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5072),
    .DIN2_t(n5072_t),
    .Q(WX9847),
    .Q_t(WX9847_t)
  );


  and2s3
  U53
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5076),
    .DIN2_t(n5076_t),
    .Q(WX9845),
    .Q_t(WX9845_t)
  );


  and2s3
  U54
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5080),
    .DIN2_t(n5080_t),
    .Q(WX9843),
    .Q_t(WX9843_t)
  );


  and2s3
  U55
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5084),
    .DIN2_t(n5084_t),
    .Q(WX9841),
    .Q_t(WX9841_t)
  );


  and2s3
  U56
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5088),
    .DIN2_t(n5088_t),
    .Q(WX9839),
    .Q_t(WX9839_t)
  );


  and2s3
  U57
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5092),
    .DIN2_t(n5092_t),
    .Q(WX9837),
    .Q_t(WX9837_t)
  );


  and2s3
  U58
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5096),
    .DIN2_t(n5096_t),
    .Q(WX9835),
    .Q_t(WX9835_t)
  );


  and2s3
  U59
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5100),
    .DIN2_t(n5100_t),
    .Q(WX9833),
    .Q_t(WX9833_t)
  );


  and2s3
  U60
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5104),
    .DIN2_t(n5104_t),
    .Q(WX9831),
    .Q_t(WX9831_t)
  );


  and2s3
  U61
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5108),
    .DIN2_t(n5108_t),
    .Q(WX9829),
    .Q_t(WX9829_t)
  );


  and2s3
  U62
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5112),
    .DIN2_t(n5112_t),
    .Q(WX9827),
    .Q_t(WX9827_t)
  );


  and2s3
  U63
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5116),
    .DIN2_t(n5116_t),
    .Q(WX9825),
    .Q_t(WX9825_t)
  );


  and2s3
  U64
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5120),
    .DIN2_t(n5120_t),
    .Q(WX9823),
    .Q_t(WX9823_t)
  );


  and2s3
  U65
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n4995),
    .DIN2_t(n4995_t),
    .Q(WX9821),
    .Q_t(WX9821_t)
  );


  and2s3
  U66
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n4999),
    .DIN2_t(n4999_t),
    .Q(WX9819),
    .Q_t(WX9819_t)
  );


  and2s3
  U67
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5003),
    .DIN2_t(n5003_t),
    .Q(WX9817),
    .Q_t(WX9817_t)
  );


  and2s3
  U68
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5007),
    .DIN2_t(n5007_t),
    .Q(WX9815),
    .Q_t(WX9815_t)
  );


  and2s3
  U69
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5011),
    .DIN2_t(n5011_t),
    .Q(WX9813),
    .Q_t(WX9813_t)
  );


  and2s3
  U70
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5015),
    .DIN2_t(n5015_t),
    .Q(WX9811),
    .Q_t(WX9811_t)
  );


  and2s3
  U71
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5019),
    .DIN2_t(n5019_t),
    .Q(WX9809),
    .Q_t(WX9809_t)
  );


  and2s3
  U72
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5023),
    .DIN2_t(n5023_t),
    .Q(WX9807),
    .Q_t(WX9807_t)
  );


  and2s3
  U73
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5027),
    .DIN2_t(n5027_t),
    .Q(WX9805),
    .Q_t(WX9805_t)
  );


  and2s3
  U74
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5031),
    .DIN2_t(n5031_t),
    .Q(WX9803),
    .Q_t(WX9803_t)
  );


  and2s3
  U75
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5035),
    .DIN2_t(n5035_t),
    .Q(WX9801),
    .Q_t(WX9801_t)
  );


  and2s3
  U76
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5039),
    .DIN2_t(n5039_t),
    .Q(WX9799),
    .Q_t(WX9799_t)
  );


  and2s3
  U77
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5043),
    .DIN2_t(n5043_t),
    .Q(WX9797),
    .Q_t(WX9797_t)
  );


  and2s3
  U78
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5047),
    .DIN2_t(n5047_t),
    .Q(WX9795),
    .Q_t(WX9795_t)
  );


  and2s3
  U79
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5051),
    .DIN2_t(n5051_t),
    .Q(WX9793),
    .Q_t(WX9793_t)
  );


  and2s3
  U80
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5055),
    .DIN2_t(n5055_t),
    .Q(WX9791),
    .Q_t(WX9791_t)
  );


  nor2s3
  U81
  (
    .DIN1(n5059),
    .DIN1_t(n5059_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9789),
    .Q_t(WX9789_t)
  );


  nor2s3
  U82
  (
    .DIN1(n5063),
    .DIN1_t(n5063_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9787),
    .Q_t(WX9787_t)
  );


  nor2s3
  U83
  (
    .DIN1(n5067),
    .DIN1_t(n5067_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9785),
    .Q_t(WX9785_t)
  );


  nor2s3
  U84
  (
    .DIN1(n5071),
    .DIN1_t(n5071_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9783),
    .Q_t(WX9783_t)
  );


  nor2s3
  U85
  (
    .DIN1(n5075),
    .DIN1_t(n5075_t),
    .DIN2(n6741),
    .DIN2_t(n6741_t),
    .Q(WX9781),
    .Q_t(WX9781_t)
  );


  nor2s3
  U86
  (
    .DIN1(n5079),
    .DIN1_t(n5079_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9779),
    .Q_t(WX9779_t)
  );


  nor2s3
  U87
  (
    .DIN1(n5083),
    .DIN1_t(n5083_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9777),
    .Q_t(WX9777_t)
  );


  nor2s3
  U88
  (
    .DIN1(n5087),
    .DIN1_t(n5087_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9775),
    .Q_t(WX9775_t)
  );


  nor2s3
  U89
  (
    .DIN1(n5091),
    .DIN1_t(n5091_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9773),
    .Q_t(WX9773_t)
  );


  nor2s3
  U90
  (
    .DIN1(n5095),
    .DIN1_t(n5095_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9771),
    .Q_t(WX9771_t)
  );


  nor2s3
  U91
  (
    .DIN1(n5099),
    .DIN1_t(n5099_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9769),
    .Q_t(WX9769_t)
  );


  nor2s3
  U92
  (
    .DIN1(n5103),
    .DIN1_t(n5103_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9767),
    .Q_t(WX9767_t)
  );


  nor2s3
  U93
  (
    .DIN1(n5107),
    .DIN1_t(n5107_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9765),
    .Q_t(WX9765_t)
  );


  nor2s3
  U94
  (
    .DIN1(n5111),
    .DIN1_t(n5111_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9763),
    .Q_t(WX9763_t)
  );


  nor2s3
  U95
  (
    .DIN1(n5115),
    .DIN1_t(n5115_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9761),
    .Q_t(WX9761_t)
  );


  nor2s3
  U96
  (
    .DIN1(n5119),
    .DIN1_t(n5119_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9759),
    .Q_t(WX9759_t)
  );


  nnd4s2
  U97
  (
    .DIN1(n2308),
    .DIN1_t(n2308_t),
    .DIN2(n2309),
    .DIN2_t(n2309_t),
    .DIN3(n2310),
    .DIN3_t(n2310_t),
    .DIN4(n2311),
    .DIN4_t(n2311_t),
    .Q(WX9757),
    .Q_t(WX9757_t)
  );


  nnd2s3
  U98
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n2313),
    .DIN2_t(n2313_t),
    .Q(n2311),
    .Q_t(n2311_t)
  );


  nnd2s3
  U99
  (
    .DIN1(n6625),
    .DIN1_t(n6625_t),
    .DIN2(n2315),
    .DIN2_t(n2315_t),
    .Q(n2310),
    .Q_t(n2310_t)
  );


  nnd2s3
  U100
  (
    .DIN1(n6616),
    .DIN1_t(n6616_t),
    .DIN2(n1825),
    .DIN2_t(n1825_t),
    .Q(n2309),
    .Q_t(n2309_t)
  );


  nnd2s3
  U101
  (
    .DIN1(n6585),
    .DIN1_t(n6585_t),
    .DIN2(n1824),
    .DIN2_t(n1824_t),
    .Q(n2308),
    .Q_t(n2308_t)
  );


  nnd4s2
  U102
  (
    .DIN1(n2318),
    .DIN1_t(n2318_t),
    .DIN2(n2319),
    .DIN2_t(n2319_t),
    .DIN3(n2320),
    .DIN3_t(n2320_t),
    .DIN4(n2321),
    .DIN4_t(n2321_t),
    .Q(WX9755),
    .Q_t(WX9755_t)
  );


  nnd2s3
  U103
  (
    .DIN1(n2322),
    .DIN1_t(n2322_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n2321),
    .Q_t(n2321_t)
  );


  nnd2s3
  U104
  (
    .DIN1(n2323),
    .DIN1_t(n2323_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n2320),
    .Q_t(n2320_t)
  );


  nnd2s3
  U105
  (
    .DIN1(n6616),
    .DIN1_t(n6616_t),
    .DIN2(n1826),
    .DIN2_t(n1826_t),
    .Q(n2319),
    .Q_t(n2319_t)
  );


  nnd2s3
  U106
  (
    .DIN1(n6585),
    .DIN1_t(n6585_t),
    .DIN2(n1823),
    .DIN2_t(n1823_t),
    .Q(n2318),
    .Q_t(n2318_t)
  );


  nnd4s2
  U107
  (
    .DIN1(n2324),
    .DIN1_t(n2324_t),
    .DIN2(n2325),
    .DIN2_t(n2325_t),
    .DIN3(n2326),
    .DIN3_t(n2326_t),
    .DIN4(n2327),
    .DIN4_t(n2327_t),
    .Q(WX9753),
    .Q_t(WX9753_t)
  );


  nnd2s3
  U108
  (
    .DIN1(n2328),
    .DIN1_t(n2328_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2327),
    .Q_t(n2327_t)
  );


  nnd2s3
  U109
  (
    .DIN1(n2329),
    .DIN1_t(n2329_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2326),
    .Q_t(n2326_t)
  );


  nnd2s3
  U110
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1827),
    .DIN2_t(n1827_t),
    .Q(n2325),
    .Q_t(n2325_t)
  );


  nnd2s3
  U111
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1822),
    .DIN2_t(n1822_t),
    .Q(n2324),
    .Q_t(n2324_t)
  );


  nnd4s2
  U112
  (
    .DIN1(n2330),
    .DIN1_t(n2330_t),
    .DIN2(n2331),
    .DIN2_t(n2331_t),
    .DIN3(n2332),
    .DIN3_t(n2332_t),
    .DIN4(n2333),
    .DIN4_t(n2333_t),
    .Q(WX9751),
    .Q_t(WX9751_t)
  );


  nnd2s3
  U113
  (
    .DIN1(n2334),
    .DIN1_t(n2334_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2333),
    .Q_t(n2333_t)
  );


  nnd2s3
  U114
  (
    .DIN1(n2335),
    .DIN1_t(n2335_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2332),
    .Q_t(n2332_t)
  );


  nnd2s3
  U115
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1828),
    .DIN2_t(n1828_t),
    .Q(n2331),
    .Q_t(n2331_t)
  );


  nnd2s3
  U116
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1821),
    .DIN2_t(n1821_t),
    .Q(n2330),
    .Q_t(n2330_t)
  );


  nnd4s2
  U117
  (
    .DIN1(n2336),
    .DIN1_t(n2336_t),
    .DIN2(n2337),
    .DIN2_t(n2337_t),
    .DIN3(n2338),
    .DIN3_t(n2338_t),
    .DIN4(n2339),
    .DIN4_t(n2339_t),
    .Q(WX9749),
    .Q_t(WX9749_t)
  );


  nnd2s3
  U118
  (
    .DIN1(n2340),
    .DIN1_t(n2340_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2339),
    .Q_t(n2339_t)
  );


  nnd2s3
  U119
  (
    .DIN1(n2341),
    .DIN1_t(n2341_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2338),
    .Q_t(n2338_t)
  );


  nnd2s3
  U120
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1829),
    .DIN2_t(n1829_t),
    .Q(n2337),
    .Q_t(n2337_t)
  );


  nnd2s3
  U121
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1820),
    .DIN2_t(n1820_t),
    .Q(n2336),
    .Q_t(n2336_t)
  );


  nnd4s2
  U122
  (
    .DIN1(n2342),
    .DIN1_t(n2342_t),
    .DIN2(n2343),
    .DIN2_t(n2343_t),
    .DIN3(n2344),
    .DIN3_t(n2344_t),
    .DIN4(n2345),
    .DIN4_t(n2345_t),
    .Q(WX9747),
    .Q_t(WX9747_t)
  );


  nnd2s3
  U123
  (
    .DIN1(n2346),
    .DIN1_t(n2346_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2345),
    .Q_t(n2345_t)
  );


  nnd2s3
  U124
  (
    .DIN1(n2347),
    .DIN1_t(n2347_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2344),
    .Q_t(n2344_t)
  );


  nnd2s3
  U125
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1830),
    .DIN2_t(n1830_t),
    .Q(n2343),
    .Q_t(n2343_t)
  );


  nnd2s3
  U126
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1819),
    .DIN2_t(n1819_t),
    .Q(n2342),
    .Q_t(n2342_t)
  );


  nnd4s2
  U127
  (
    .DIN1(n2348),
    .DIN1_t(n2348_t),
    .DIN2(n2349),
    .DIN2_t(n2349_t),
    .DIN3(n2350),
    .DIN3_t(n2350_t),
    .DIN4(n2351),
    .DIN4_t(n2351_t),
    .Q(WX9745),
    .Q_t(WX9745_t)
  );


  nnd2s3
  U128
  (
    .DIN1(n2352),
    .DIN1_t(n2352_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2351),
    .Q_t(n2351_t)
  );


  nnd2s3
  U129
  (
    .DIN1(n2353),
    .DIN1_t(n2353_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2350),
    .Q_t(n2350_t)
  );


  nnd2s3
  U130
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1831),
    .DIN2_t(n1831_t),
    .Q(n2349),
    .Q_t(n2349_t)
  );


  nnd2s3
  U131
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1818),
    .DIN2_t(n1818_t),
    .Q(n2348),
    .Q_t(n2348_t)
  );


  nnd4s2
  U132
  (
    .DIN1(n2354),
    .DIN1_t(n2354_t),
    .DIN2(n2355),
    .DIN2_t(n2355_t),
    .DIN3(n2356),
    .DIN3_t(n2356_t),
    .DIN4(n2357),
    .DIN4_t(n2357_t),
    .Q(WX9743),
    .Q_t(WX9743_t)
  );


  nnd2s3
  U133
  (
    .DIN1(n2358),
    .DIN1_t(n2358_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2357),
    .Q_t(n2357_t)
  );


  nnd2s3
  U134
  (
    .DIN1(n2359),
    .DIN1_t(n2359_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2356),
    .Q_t(n2356_t)
  );


  nnd2s3
  U135
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1832),
    .DIN2_t(n1832_t),
    .Q(n2355),
    .Q_t(n2355_t)
  );


  nnd2s3
  U136
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1817),
    .DIN2_t(n1817_t),
    .Q(n2354),
    .Q_t(n2354_t)
  );


  nnd4s2
  U137
  (
    .DIN1(n2360),
    .DIN1_t(n2360_t),
    .DIN2(n2361),
    .DIN2_t(n2361_t),
    .DIN3(n2362),
    .DIN3_t(n2362_t),
    .DIN4(n2363),
    .DIN4_t(n2363_t),
    .Q(WX9741),
    .Q_t(WX9741_t)
  );


  nnd2s3
  U138
  (
    .DIN1(n2364),
    .DIN1_t(n2364_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2363),
    .Q_t(n2363_t)
  );


  nnd2s3
  U139
  (
    .DIN1(n2365),
    .DIN1_t(n2365_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2362),
    .Q_t(n2362_t)
  );


  nnd2s3
  U140
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1833),
    .DIN2_t(n1833_t),
    .Q(n2361),
    .Q_t(n2361_t)
  );


  nnd2s3
  U141
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1816),
    .DIN2_t(n1816_t),
    .Q(n2360),
    .Q_t(n2360_t)
  );


  nnd4s2
  U142
  (
    .DIN1(n2366),
    .DIN1_t(n2366_t),
    .DIN2(n2367),
    .DIN2_t(n2367_t),
    .DIN3(n2368),
    .DIN3_t(n2368_t),
    .DIN4(n2369),
    .DIN4_t(n2369_t),
    .Q(WX9739),
    .Q_t(WX9739_t)
  );


  nnd2s3
  U143
  (
    .DIN1(n2370),
    .DIN1_t(n2370_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2369),
    .Q_t(n2369_t)
  );


  nnd2s3
  U144
  (
    .DIN1(n2371),
    .DIN1_t(n2371_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2368),
    .Q_t(n2368_t)
  );


  nnd2s3
  U145
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1834),
    .DIN2_t(n1834_t),
    .Q(n2367),
    .Q_t(n2367_t)
  );


  nnd2s3
  U146
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1815),
    .DIN2_t(n1815_t),
    .Q(n2366),
    .Q_t(n2366_t)
  );


  nnd4s2
  U147
  (
    .DIN1(n2372),
    .DIN1_t(n2372_t),
    .DIN2(n2373),
    .DIN2_t(n2373_t),
    .DIN3(n2374),
    .DIN3_t(n2374_t),
    .DIN4(n2375),
    .DIN4_t(n2375_t),
    .Q(WX9737),
    .Q_t(WX9737_t)
  );


  nnd2s3
  U148
  (
    .DIN1(n2376),
    .DIN1_t(n2376_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2375),
    .Q_t(n2375_t)
  );


  nnd2s3
  U149
  (
    .DIN1(n2377),
    .DIN1_t(n2377_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2374),
    .Q_t(n2374_t)
  );


  nnd2s3
  U150
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1835),
    .DIN2_t(n1835_t),
    .Q(n2373),
    .Q_t(n2373_t)
  );


  nnd2s3
  U151
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1814),
    .DIN2_t(n1814_t),
    .Q(n2372),
    .Q_t(n2372_t)
  );


  nnd4s2
  U152
  (
    .DIN1(n2378),
    .DIN1_t(n2378_t),
    .DIN2(n2379),
    .DIN2_t(n2379_t),
    .DIN3(n2380),
    .DIN3_t(n2380_t),
    .DIN4(n2381),
    .DIN4_t(n2381_t),
    .Q(WX9735),
    .Q_t(WX9735_t)
  );


  nnd2s3
  U153
  (
    .DIN1(n2382),
    .DIN1_t(n2382_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2381),
    .Q_t(n2381_t)
  );


  nnd2s3
  U154
  (
    .DIN1(n2383),
    .DIN1_t(n2383_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2380),
    .Q_t(n2380_t)
  );


  nnd2s3
  U155
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1836),
    .DIN2_t(n1836_t),
    .Q(n2379),
    .Q_t(n2379_t)
  );


  nnd2s3
  U156
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1813),
    .DIN2_t(n1813_t),
    .Q(n2378),
    .Q_t(n2378_t)
  );


  nnd4s2
  U157
  (
    .DIN1(n2384),
    .DIN1_t(n2384_t),
    .DIN2(n2385),
    .DIN2_t(n2385_t),
    .DIN3(n2386),
    .DIN3_t(n2386_t),
    .DIN4(n2387),
    .DIN4_t(n2387_t),
    .Q(WX9733),
    .Q_t(WX9733_t)
  );


  nnd2s3
  U158
  (
    .DIN1(n2388),
    .DIN1_t(n2388_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2387),
    .Q_t(n2387_t)
  );


  nnd2s3
  U159
  (
    .DIN1(n2389),
    .DIN1_t(n2389_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2386),
    .Q_t(n2386_t)
  );


  nnd2s3
  U160
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1837),
    .DIN2_t(n1837_t),
    .Q(n2385),
    .Q_t(n2385_t)
  );


  nnd2s3
  U161
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1812),
    .DIN2_t(n1812_t),
    .Q(n2384),
    .Q_t(n2384_t)
  );


  nnd4s2
  U162
  (
    .DIN1(n2390),
    .DIN1_t(n2390_t),
    .DIN2(n2391),
    .DIN2_t(n2391_t),
    .DIN3(n2392),
    .DIN3_t(n2392_t),
    .DIN4(n2393),
    .DIN4_t(n2393_t),
    .Q(WX9731),
    .Q_t(WX9731_t)
  );


  nnd2s3
  U163
  (
    .DIN1(n2394),
    .DIN1_t(n2394_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2393),
    .Q_t(n2393_t)
  );


  nnd2s3
  U164
  (
    .DIN1(n2395),
    .DIN1_t(n2395_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2392),
    .Q_t(n2392_t)
  );


  nnd2s3
  U165
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1838),
    .DIN2_t(n1838_t),
    .Q(n2391),
    .Q_t(n2391_t)
  );


  nnd2s3
  U166
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1811),
    .DIN2_t(n1811_t),
    .Q(n2390),
    .Q_t(n2390_t)
  );


  nnd4s2
  U167
  (
    .DIN1(n2396),
    .DIN1_t(n2396_t),
    .DIN2(n2397),
    .DIN2_t(n2397_t),
    .DIN3(n2398),
    .DIN3_t(n2398_t),
    .DIN4(n2399),
    .DIN4_t(n2399_t),
    .Q(WX9729),
    .Q_t(WX9729_t)
  );


  nnd2s3
  U168
  (
    .DIN1(n2400),
    .DIN1_t(n2400_t),
    .DIN2(n6666),
    .DIN2_t(n6666_t),
    .Q(n2399),
    .Q_t(n2399_t)
  );


  nnd2s3
  U169
  (
    .DIN1(n2401),
    .DIN1_t(n2401_t),
    .DIN2(n6635),
    .DIN2_t(n6635_t),
    .Q(n2398),
    .Q_t(n2398_t)
  );


  nnd2s3
  U170
  (
    .DIN1(n6615),
    .DIN1_t(n6615_t),
    .DIN2(n1839),
    .DIN2_t(n1839_t),
    .Q(n2397),
    .Q_t(n2397_t)
  );


  nnd2s3
  U171
  (
    .DIN1(n6584),
    .DIN1_t(n6584_t),
    .DIN2(n1810),
    .DIN2_t(n1810_t),
    .Q(n2396),
    .Q_t(n2396_t)
  );


  nnd4s2
  U172
  (
    .DIN1(n2402),
    .DIN1_t(n2402_t),
    .DIN2(n2403),
    .DIN2_t(n2403_t),
    .DIN3(n2404),
    .DIN3_t(n2404_t),
    .DIN4(n2405),
    .DIN4_t(n2405_t),
    .Q(WX9727),
    .Q_t(WX9727_t)
  );


  nnd2s3
  U173
  (
    .DIN1(n2406),
    .DIN1_t(n2406_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2405),
    .Q_t(n2405_t)
  );


  nnd2s3
  U174
  (
    .DIN1(n2407),
    .DIN1_t(n2407_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2404),
    .Q_t(n2404_t)
  );


  nnd2s3
  U175
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1840),
    .DIN2_t(n1840_t),
    .Q(n2403),
    .Q_t(n2403_t)
  );


  nnd2s3
  U176
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1809),
    .DIN2_t(n1809_t),
    .Q(n2402),
    .Q_t(n2402_t)
  );


  nnd4s2
  U177
  (
    .DIN1(n2408),
    .DIN1_t(n2408_t),
    .DIN2(n2409),
    .DIN2_t(n2409_t),
    .DIN3(n2410),
    .DIN3_t(n2410_t),
    .DIN4(n2411),
    .DIN4_t(n2411_t),
    .Q(WX9725),
    .Q_t(WX9725_t)
  );


  nnd2s3
  U178
  (
    .DIN1(n2412),
    .DIN1_t(n2412_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2411),
    .Q_t(n2411_t)
  );


  nnd2s3
  U179
  (
    .DIN1(n2413),
    .DIN1_t(n2413_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2410),
    .Q_t(n2410_t)
  );


  nnd2s3
  U180
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1841),
    .DIN2_t(n1841_t),
    .Q(n2409),
    .Q_t(n2409_t)
  );


  nnd2s3
  U181
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1808),
    .DIN2_t(n1808_t),
    .Q(n2408),
    .Q_t(n2408_t)
  );


  nnd4s2
  U182
  (
    .DIN1(n2414),
    .DIN1_t(n2414_t),
    .DIN2(n2415),
    .DIN2_t(n2415_t),
    .DIN3(n2416),
    .DIN3_t(n2416_t),
    .DIN4(n2417),
    .DIN4_t(n2417_t),
    .Q(WX9723),
    .Q_t(WX9723_t)
  );


  nnd2s3
  U183
  (
    .DIN1(n2418),
    .DIN1_t(n2418_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2417),
    .Q_t(n2417_t)
  );


  nnd2s3
  U184
  (
    .DIN1(n2419),
    .DIN1_t(n2419_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2416),
    .Q_t(n2416_t)
  );


  nnd2s3
  U185
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1842),
    .DIN2_t(n1842_t),
    .Q(n2415),
    .Q_t(n2415_t)
  );


  nnd2s3
  U186
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1807),
    .DIN2_t(n1807_t),
    .Q(n2414),
    .Q_t(n2414_t)
  );


  nnd4s2
  U187
  (
    .DIN1(n2420),
    .DIN1_t(n2420_t),
    .DIN2(n2421),
    .DIN2_t(n2421_t),
    .DIN3(n2422),
    .DIN3_t(n2422_t),
    .DIN4(n2423),
    .DIN4_t(n2423_t),
    .Q(WX9721),
    .Q_t(WX9721_t)
  );


  nnd2s3
  U188
  (
    .DIN1(n2424),
    .DIN1_t(n2424_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2423),
    .Q_t(n2423_t)
  );


  nnd2s3
  U189
  (
    .DIN1(n2425),
    .DIN1_t(n2425_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2422),
    .Q_t(n2422_t)
  );


  nnd2s3
  U190
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1843),
    .DIN2_t(n1843_t),
    .Q(n2421),
    .Q_t(n2421_t)
  );


  nnd2s3
  U191
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1806),
    .DIN2_t(n1806_t),
    .Q(n2420),
    .Q_t(n2420_t)
  );


  nnd4s2
  U192
  (
    .DIN1(n2426),
    .DIN1_t(n2426_t),
    .DIN2(n2427),
    .DIN2_t(n2427_t),
    .DIN3(n2428),
    .DIN3_t(n2428_t),
    .DIN4(n2429),
    .DIN4_t(n2429_t),
    .Q(WX9719),
    .Q_t(WX9719_t)
  );


  nnd2s3
  U193
  (
    .DIN1(n2430),
    .DIN1_t(n2430_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2429),
    .Q_t(n2429_t)
  );


  nnd2s3
  U194
  (
    .DIN1(n2431),
    .DIN1_t(n2431_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2428),
    .Q_t(n2428_t)
  );


  nnd2s3
  U195
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1844),
    .DIN2_t(n1844_t),
    .Q(n2427),
    .Q_t(n2427_t)
  );


  nnd2s3
  U196
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1805),
    .DIN2_t(n1805_t),
    .Q(n2426),
    .Q_t(n2426_t)
  );


  nnd4s2
  U197
  (
    .DIN1(n2432),
    .DIN1_t(n2432_t),
    .DIN2(n2433),
    .DIN2_t(n2433_t),
    .DIN3(n2434),
    .DIN3_t(n2434_t),
    .DIN4(n2435),
    .DIN4_t(n2435_t),
    .Q(WX9717),
    .Q_t(WX9717_t)
  );


  nnd2s3
  U198
  (
    .DIN1(n2436),
    .DIN1_t(n2436_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2435),
    .Q_t(n2435_t)
  );


  nnd2s3
  U199
  (
    .DIN1(n2437),
    .DIN1_t(n2437_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2434),
    .Q_t(n2434_t)
  );


  nnd2s3
  U200
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1845),
    .DIN2_t(n1845_t),
    .Q(n2433),
    .Q_t(n2433_t)
  );


  nnd2s3
  U201
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1804),
    .DIN2_t(n1804_t),
    .Q(n2432),
    .Q_t(n2432_t)
  );


  nnd4s2
  U202
  (
    .DIN1(n2438),
    .DIN1_t(n2438_t),
    .DIN2(n2439),
    .DIN2_t(n2439_t),
    .DIN3(n2440),
    .DIN3_t(n2440_t),
    .DIN4(n2441),
    .DIN4_t(n2441_t),
    .Q(WX9715),
    .Q_t(WX9715_t)
  );


  nnd2s3
  U203
  (
    .DIN1(n2442),
    .DIN1_t(n2442_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2441),
    .Q_t(n2441_t)
  );


  nnd2s3
  U204
  (
    .DIN1(n2443),
    .DIN1_t(n2443_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2440),
    .Q_t(n2440_t)
  );


  nnd2s3
  U205
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1846),
    .DIN2_t(n1846_t),
    .Q(n2439),
    .Q_t(n2439_t)
  );


  nnd2s3
  U206
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1803),
    .DIN2_t(n1803_t),
    .Q(n2438),
    .Q_t(n2438_t)
  );


  nnd4s2
  U207
  (
    .DIN1(n2444),
    .DIN1_t(n2444_t),
    .DIN2(n2445),
    .DIN2_t(n2445_t),
    .DIN3(n2446),
    .DIN3_t(n2446_t),
    .DIN4(n2447),
    .DIN4_t(n2447_t),
    .Q(WX9713),
    .Q_t(WX9713_t)
  );


  nnd2s3
  U208
  (
    .DIN1(n2448),
    .DIN1_t(n2448_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2447),
    .Q_t(n2447_t)
  );


  nnd2s3
  U209
  (
    .DIN1(n2449),
    .DIN1_t(n2449_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2446),
    .Q_t(n2446_t)
  );


  nnd2s3
  U210
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1847),
    .DIN2_t(n1847_t),
    .Q(n2445),
    .Q_t(n2445_t)
  );


  nnd2s3
  U211
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1802),
    .DIN2_t(n1802_t),
    .Q(n2444),
    .Q_t(n2444_t)
  );


  nnd4s2
  U212
  (
    .DIN1(n2450),
    .DIN1_t(n2450_t),
    .DIN2(n2451),
    .DIN2_t(n2451_t),
    .DIN3(n2452),
    .DIN3_t(n2452_t),
    .DIN4(n2453),
    .DIN4_t(n2453_t),
    .Q(WX9711),
    .Q_t(WX9711_t)
  );


  nnd2s3
  U213
  (
    .DIN1(n2454),
    .DIN1_t(n2454_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2453),
    .Q_t(n2453_t)
  );


  nnd2s3
  U214
  (
    .DIN1(n2455),
    .DIN1_t(n2455_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2452),
    .Q_t(n2452_t)
  );


  nnd2s3
  U215
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1848),
    .DIN2_t(n1848_t),
    .Q(n2451),
    .Q_t(n2451_t)
  );


  nnd2s3
  U216
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1801),
    .DIN2_t(n1801_t),
    .Q(n2450),
    .Q_t(n2450_t)
  );


  nnd4s2
  U217
  (
    .DIN1(n2456),
    .DIN1_t(n2456_t),
    .DIN2(n2457),
    .DIN2_t(n2457_t),
    .DIN3(n2458),
    .DIN3_t(n2458_t),
    .DIN4(n2459),
    .DIN4_t(n2459_t),
    .Q(WX9709),
    .Q_t(WX9709_t)
  );


  nnd2s3
  U218
  (
    .DIN1(n2460),
    .DIN1_t(n2460_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2459),
    .Q_t(n2459_t)
  );


  nnd2s3
  U219
  (
    .DIN1(n2461),
    .DIN1_t(n2461_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2458),
    .Q_t(n2458_t)
  );


  nnd2s3
  U220
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1849),
    .DIN2_t(n1849_t),
    .Q(n2457),
    .Q_t(n2457_t)
  );


  nnd2s3
  U221
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1800),
    .DIN2_t(n1800_t),
    .Q(n2456),
    .Q_t(n2456_t)
  );


  nnd4s2
  U222
  (
    .DIN1(n2462),
    .DIN1_t(n2462_t),
    .DIN2(n2463),
    .DIN2_t(n2463_t),
    .DIN3(n2464),
    .DIN3_t(n2464_t),
    .DIN4(n2465),
    .DIN4_t(n2465_t),
    .Q(WX9707),
    .Q_t(WX9707_t)
  );


  nnd2s3
  U223
  (
    .DIN1(n2466),
    .DIN1_t(n2466_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2465),
    .Q_t(n2465_t)
  );


  nnd2s3
  U224
  (
    .DIN1(n2467),
    .DIN1_t(n2467_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2464),
    .Q_t(n2464_t)
  );


  nnd2s3
  U225
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1850),
    .DIN2_t(n1850_t),
    .Q(n2463),
    .Q_t(n2463_t)
  );


  nnd2s3
  U226
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1799),
    .DIN2_t(n1799_t),
    .Q(n2462),
    .Q_t(n2462_t)
  );


  nnd4s2
  U227
  (
    .DIN1(n2468),
    .DIN1_t(n2468_t),
    .DIN2(n2469),
    .DIN2_t(n2469_t),
    .DIN3(n2470),
    .DIN3_t(n2470_t),
    .DIN4(n2471),
    .DIN4_t(n2471_t),
    .Q(WX9705),
    .Q_t(WX9705_t)
  );


  nnd2s3
  U228
  (
    .DIN1(n2472),
    .DIN1_t(n2472_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2471),
    .Q_t(n2471_t)
  );


  nnd2s3
  U229
  (
    .DIN1(n2473),
    .DIN1_t(n2473_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2470),
    .Q_t(n2470_t)
  );


  nnd2s3
  U230
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1851),
    .DIN2_t(n1851_t),
    .Q(n2469),
    .Q_t(n2469_t)
  );


  nnd2s3
  U231
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1798),
    .DIN2_t(n1798_t),
    .Q(n2468),
    .Q_t(n2468_t)
  );


  nnd4s2
  U232
  (
    .DIN1(n2474),
    .DIN1_t(n2474_t),
    .DIN2(n2475),
    .DIN2_t(n2475_t),
    .DIN3(n2476),
    .DIN3_t(n2476_t),
    .DIN4(n2477),
    .DIN4_t(n2477_t),
    .Q(WX9703),
    .Q_t(WX9703_t)
  );


  nnd2s3
  U233
  (
    .DIN1(n2478),
    .DIN1_t(n2478_t),
    .DIN2(n6665),
    .DIN2_t(n6665_t),
    .Q(n2477),
    .Q_t(n2477_t)
  );


  nnd2s3
  U234
  (
    .DIN1(n2479),
    .DIN1_t(n2479_t),
    .DIN2(n6634),
    .DIN2_t(n6634_t),
    .Q(n2476),
    .Q_t(n2476_t)
  );


  nnd2s3
  U235
  (
    .DIN1(n6614),
    .DIN1_t(n6614_t),
    .DIN2(n1852),
    .DIN2_t(n1852_t),
    .Q(n2475),
    .Q_t(n2475_t)
  );


  nnd2s3
  U236
  (
    .DIN1(n6583),
    .DIN1_t(n6583_t),
    .DIN2(n1797),
    .DIN2_t(n1797_t),
    .Q(n2474),
    .Q_t(n2474_t)
  );


  nnd4s2
  U237
  (
    .DIN1(n2480),
    .DIN1_t(n2480_t),
    .DIN2(n2481),
    .DIN2_t(n2481_t),
    .DIN3(n2482),
    .DIN3_t(n2482_t),
    .DIN4(n2483),
    .DIN4_t(n2483_t),
    .Q(WX9701),
    .Q_t(WX9701_t)
  );


  nnd2s3
  U238
  (
    .DIN1(n2484),
    .DIN1_t(n2484_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2483),
    .Q_t(n2483_t)
  );


  nnd2s3
  U239
  (
    .DIN1(n2485),
    .DIN1_t(n2485_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2482),
    .Q_t(n2482_t)
  );


  nnd2s3
  U240
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1853),
    .DIN2_t(n1853_t),
    .Q(n2481),
    .Q_t(n2481_t)
  );


  nnd2s3
  U241
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1796),
    .DIN2_t(n1796_t),
    .Q(n2480),
    .Q_t(n2480_t)
  );


  nnd4s2
  U242
  (
    .DIN1(n2486),
    .DIN1_t(n2486_t),
    .DIN2(n2487),
    .DIN2_t(n2487_t),
    .DIN3(n2488),
    .DIN3_t(n2488_t),
    .DIN4(n2489),
    .DIN4_t(n2489_t),
    .Q(WX9699),
    .Q_t(WX9699_t)
  );


  nnd2s3
  U243
  (
    .DIN1(n2490),
    .DIN1_t(n2490_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2489),
    .Q_t(n2489_t)
  );


  nnd2s3
  U244
  (
    .DIN1(n2491),
    .DIN1_t(n2491_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2488),
    .Q_t(n2488_t)
  );


  nnd2s3
  U245
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1854),
    .DIN2_t(n1854_t),
    .Q(n2487),
    .Q_t(n2487_t)
  );


  nnd2s3
  U246
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1795),
    .DIN2_t(n1795_t),
    .Q(n2486),
    .Q_t(n2486_t)
  );


  nnd4s2
  U247
  (
    .DIN1(n2492),
    .DIN1_t(n2492_t),
    .DIN2(n2493),
    .DIN2_t(n2493_t),
    .DIN3(n2494),
    .DIN3_t(n2494_t),
    .DIN4(n2495),
    .DIN4_t(n2495_t),
    .Q(WX9697),
    .Q_t(WX9697_t)
  );


  nnd2s3
  U248
  (
    .DIN1(n2496),
    .DIN1_t(n2496_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2495),
    .Q_t(n2495_t)
  );


  nnd2s3
  U249
  (
    .DIN1(n2497),
    .DIN1_t(n2497_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2494),
    .Q_t(n2494_t)
  );


  nnd2s3
  U250
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1855),
    .DIN2_t(n1855_t),
    .Q(tempn2493),
    .Q_t(tempn2493_t)
  );


  nnd2s3
  U251
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1794),
    .DIN2_t(n1794_t),
    .Q(n2492),
    .Q_t(n2492_t)
  );


  nnd4s2
  U252
  (
    .DIN1(n2498),
    .DIN1_t(n2498_t),
    .DIN2(n2499),
    .DIN2_t(n2499_t),
    .DIN3(n2500),
    .DIN3_t(n2500_t),
    .DIN4(n2501),
    .DIN4_t(n2501_t),
    .Q(WX9695),
    .Q_t(WX9695_t)
  );


  nnd2s3
  U253
  (
    .DIN1(n2502),
    .DIN1_t(n2502_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2501),
    .Q_t(n2501_t)
  );


  nnd2s3
  U254
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1856),
    .DIN2_t(n1856_t),
    .Q(n2500),
    .Q_t(n2500_t)
  );


  nnd2s3
  U255
  (
    .DIN1(n2503),
    .DIN1_t(n2503_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2499),
    .Q_t(n2499_t)
  );


  nnd2s3
  U256
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1793),
    .DIN2_t(n1793_t),
    .Q(n2498),
    .Q_t(n2498_t)
  );


  nor2s3
  U257
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n1856),
    .DIN2_t(n1856_t),
    .Q(WX9597),
    .Q_t(WX9597_t)
  );


  nor2s3
  U258
  (
    .DIN1(n4964),
    .DIN1_t(n4964_t),
    .DIN2(n6740),
    .DIN2_t(n6740_t),
    .Q(WX9595),
    .Q_t(WX9595_t)
  );


  nor2s3
  U259
  (
    .DIN1(n4965),
    .DIN1_t(n4965_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX9593),
    .Q_t(WX9593_t)
  );


  nor2s3
  U260
  (
    .DIN1(n4966),
    .DIN1_t(n4966_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX9591),
    .Q_t(WX9591_t)
  );


  nor2s3
  U261
  (
    .DIN1(n4967),
    .DIN1_t(n4967_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX9589),
    .Q_t(WX9589_t)
  );


  nor2s3
  U262
  (
    .DIN1(n4968),
    .DIN1_t(n4968_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX9587),
    .Q_t(WX9587_t)
  );


  nor2s3
  U263
  (
    .DIN1(n4969),
    .DIN1_t(n4969_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX9585),
    .Q_t(WX9585_t)
  );


  nor2s3
  U264
  (
    .DIN1(n4970),
    .DIN1_t(n4970_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX9583),
    .Q_t(WX9583_t)
  );


  nor2s3
  U265
  (
    .DIN1(n4971),
    .DIN1_t(n4971_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX9581),
    .Q_t(WX9581_t)
  );


  nor2s3
  U266
  (
    .DIN1(n4972),
    .DIN1_t(n4972_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX9579),
    .Q_t(WX9579_t)
  );


  nor2s3
  U267
  (
    .DIN1(n4973),
    .DIN1_t(n4973_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX9577),
    .Q_t(WX9577_t)
  );


  nor2s3
  U268
  (
    .DIN1(n4974),
    .DIN1_t(n4974_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX9575),
    .Q_t(WX9575_t)
  );


  nor2s3
  U269
  (
    .DIN1(n4975),
    .DIN1_t(n4975_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX9573),
    .Q_t(WX9573_t)
  );


  nor2s3
  U270
  (
    .DIN1(n4976),
    .DIN1_t(n4976_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9571),
    .Q_t(WX9571_t)
  );


  nor2s3
  U271
  (
    .DIN1(n4977),
    .DIN1_t(n4977_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9569),
    .Q_t(WX9569_t)
  );


  nor2s3
  U272
  (
    .DIN1(n4978),
    .DIN1_t(n4978_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9567),
    .Q_t(WX9567_t)
  );


  nor2s3
  U273
  (
    .DIN1(n4979),
    .DIN1_t(n4979_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9565),
    .Q_t(WX9565_t)
  );


  nor2s3
  U274
  (
    .DIN1(n4980),
    .DIN1_t(n4980_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9563),
    .Q_t(WX9563_t)
  );


  nor2s3
  U275
  (
    .DIN1(n4981),
    .DIN1_t(n4981_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9561),
    .Q_t(WX9561_t)
  );


  nor2s3
  U276
  (
    .DIN1(n4982),
    .DIN1_t(n4982_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9559),
    .Q_t(WX9559_t)
  );


  nor2s3
  U277
  (
    .DIN1(n4983),
    .DIN1_t(n4983_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9557),
    .Q_t(WX9557_t)
  );


  nor2s3
  U278
  (
    .DIN1(n4984),
    .DIN1_t(n4984_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9555),
    .Q_t(WX9555_t)
  );


  nor2s3
  U279
  (
    .DIN1(n4985),
    .DIN1_t(n4985_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9553),
    .Q_t(WX9553_t)
  );


  nor2s3
  U280
  (
    .DIN1(n4986),
    .DIN1_t(n4986_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9551),
    .Q_t(WX9551_t)
  );


  nor2s3
  U281
  (
    .DIN1(n4987),
    .DIN1_t(n4987_t),
    .DIN2(n6738),
    .DIN2_t(n6738_t),
    .Q(WX9549),
    .Q_t(WX9549_t)
  );


  nor2s3
  U282
  (
    .DIN1(n4988),
    .DIN1_t(n4988_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX9547),
    .Q_t(WX9547_t)
  );


  nor2s3
  U283
  (
    .DIN1(n4989),
    .DIN1_t(n4989_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX9545),
    .Q_t(WX9545_t)
  );


  nor2s3
  U284
  (
    .DIN1(n4990),
    .DIN1_t(n4990_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX9543),
    .Q_t(WX9543_t)
  );


  nor2s3
  U285
  (
    .DIN1(n4991),
    .DIN1_t(n4991_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX9541),
    .Q_t(WX9541_t)
  );


  nor2s3
  U286
  (
    .DIN1(n4992),
    .DIN1_t(n4992_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX9539),
    .Q_t(WX9539_t)
  );


  nor2s3
  U287
  (
    .DIN1(n4993),
    .DIN1_t(n4993_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX9537),
    .Q_t(WX9537_t)
  );


  nor2s3
  U288
  (
    .DIN1(n4994),
    .DIN1_t(n4994_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX9535),
    .Q_t(WX9535_t)
  );


  nor2s3
  U289
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n2504),
    .DIN2_t(n2504_t),
    .Q(WX9084),
    .Q_t(WX9084_t)
  );


  xor2s3
  U290
  (
    .DIN1(n5118),
    .DIN1_t(n5118_t),
    .DIN2(n5297),
    .DIN2_t(n5297_t),
    .Q(n2504),
    .Q_t(n2504_t)
  );


  nor2s3
  U291
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n2505),
    .DIN2_t(n2505_t),
    .Q(WX9082),
    .Q_t(WX9082_t)
  );


  xor2s3
  U292
  (
    .DIN1(n5114),
    .DIN1_t(n5114_t),
    .DIN2(n5292),
    .DIN2_t(n5292_t),
    .Q(n2505),
    .Q_t(n2505_t)
  );


  nor2s3
  U293
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n2506),
    .DIN2_t(n2506_t),
    .Q(WX9080),
    .Q_t(WX9080_t)
  );


  xor2s3
  U294
  (
    .DIN1(n5110),
    .DIN1_t(n5110_t),
    .DIN2(n5287),
    .DIN2_t(n5287_t),
    .Q(n2506),
    .Q_t(n2506_t)
  );


  nor2s3
  U295
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n2507),
    .DIN2_t(n2507_t),
    .Q(WX9078),
    .Q_t(WX9078_t)
  );


  xor2s3
  U296
  (
    .DIN1(n5106),
    .DIN1_t(n5106_t),
    .DIN2(n5282),
    .DIN2_t(n5282_t),
    .Q(n2507),
    .Q_t(n2507_t)
  );


  nor2s3
  U297
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n2508),
    .DIN2_t(n2508_t),
    .Q(WX9076),
    .Q_t(WX9076_t)
  );


  xor2s3
  U298
  (
    .DIN1(n5102),
    .DIN1_t(n5102_t),
    .DIN2(n5277),
    .DIN2_t(n5277_t),
    .Q(n2508),
    .Q_t(n2508_t)
  );


  nor2s3
  U299
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n2509),
    .DIN2_t(n2509_t),
    .Q(WX9074),
    .Q_t(WX9074_t)
  );


  xor2s3
  U300
  (
    .DIN1(n5098),
    .DIN1_t(n5098_t),
    .DIN2(n5272),
    .DIN2_t(n5272_t),
    .Q(n2509),
    .Q_t(n2509_t)
  );


  nor2s3
  U301
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n2510),
    .DIN2_t(n2510_t),
    .Q(WX9072),
    .Q_t(WX9072_t)
  );


  xor2s3
  U302
  (
    .DIN1(n5094),
    .DIN1_t(n5094_t),
    .DIN2(n5267),
    .DIN2_t(n5267_t),
    .Q(n2510),
    .Q_t(n2510_t)
  );


  nor2s3
  U303
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n2511),
    .DIN2_t(n2511_t),
    .Q(WX9070),
    .Q_t(WX9070_t)
  );


  xor2s3
  U304
  (
    .DIN1(n5090),
    .DIN1_t(n5090_t),
    .DIN2(n5262),
    .DIN2_t(n5262_t),
    .Q(n2511),
    .Q_t(n2511_t)
  );


  nor2s3
  U305
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n2512),
    .DIN2_t(n2512_t),
    .Q(WX9068),
    .Q_t(WX9068_t)
  );


  xor2s3
  U306
  (
    .DIN1(n5086),
    .DIN1_t(n5086_t),
    .DIN2(n5257),
    .DIN2_t(n5257_t),
    .Q(n2512),
    .Q_t(n2512_t)
  );


  nor2s3
  U307
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n2513),
    .DIN2_t(n2513_t),
    .Q(WX9066),
    .Q_t(WX9066_t)
  );


  xor2s3
  U308
  (
    .DIN1(n5082),
    .DIN1_t(n5082_t),
    .DIN2(n5252),
    .DIN2_t(n5252_t),
    .Q(n2513),
    .Q_t(n2513_t)
  );


  nor2s3
  U309
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n2514),
    .DIN2_t(n2514_t),
    .Q(WX9064),
    .Q_t(WX9064_t)
  );


  xor2s3
  U310
  (
    .DIN1(n5078),
    .DIN1_t(n5078_t),
    .DIN2(n5247),
    .DIN2_t(n5247_t),
    .Q(n2514),
    .Q_t(n2514_t)
  );


  nor2s3
  U311
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n2515),
    .DIN2_t(n2515_t),
    .Q(WX9062),
    .Q_t(WX9062_t)
  );


  xor2s3
  U312
  (
    .DIN1(n5074),
    .DIN1_t(n5074_t),
    .DIN2(n5242),
    .DIN2_t(n5242_t),
    .Q(n2515),
    .Q_t(n2515_t)
  );


  nor2s3
  U313
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n2516),
    .DIN2_t(n2516_t),
    .Q(WX9060),
    .Q_t(WX9060_t)
  );


  xor2s3
  U314
  (
    .DIN1(n5070),
    .DIN1_t(n5070_t),
    .DIN2(n5237),
    .DIN2_t(n5237_t),
    .Q(n2516),
    .Q_t(n2516_t)
  );


  nor2s3
  U315
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n2517),
    .DIN2_t(n2517_t),
    .Q(WX9058),
    .Q_t(WX9058_t)
  );


  xor2s3
  U316
  (
    .DIN1(n5066),
    .DIN1_t(n5066_t),
    .DIN2(n5232),
    .DIN2_t(n5232_t),
    .Q(n2517),
    .Q_t(n2517_t)
  );


  nor2s3
  U317
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n2518),
    .DIN2_t(n2518_t),
    .Q(WX9056),
    .Q_t(WX9056_t)
  );


  xor2s3
  U318
  (
    .DIN1(n5062),
    .DIN1_t(n5062_t),
    .DIN2(n5227),
    .DIN2_t(n5227_t),
    .Q(n2518),
    .Q_t(n2518_t)
  );


  nor2s3
  U319
  (
    .DIN1(n2519),
    .DIN1_t(n2519_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX9054),
    .Q_t(WX9054_t)
  );


  xnr2s3
  U320
  (
    .DIN1(n5222),
    .DIN1_t(n5222_t),
    .DIN2(n2520),
    .DIN2_t(n2520_t),
    .Q(n2519),
    .Q_t(n2519_t)
  );


  xor2s3
  U321
  (
    .DIN1(n5058),
    .DIN1_t(n5058_t),
    .DIN2(n5122),
    .DIN2_t(n5122_t),
    .Q(n2520),
    .Q_t(n2520_t)
  );


  nor2s3
  U322
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n2521),
    .DIN2_t(n2521_t),
    .Q(WX9052),
    .Q_t(WX9052_t)
  );


  xor2s3
  U323
  (
    .DIN1(n5054),
    .DIN1_t(n5054_t),
    .DIN2(n3236),
    .DIN2_t(n3236_t),
    .Q(n2521),
    .Q_t(n2521_t)
  );


  nor2s3
  U324
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n2522),
    .DIN2_t(n2522_t),
    .Q(WX9050),
    .Q_t(WX9050_t)
  );


  xor2s3
  U325
  (
    .DIN1(n5050),
    .DIN1_t(n5050_t),
    .DIN2(n3235),
    .DIN2_t(n3235_t),
    .Q(n2522),
    .Q_t(n2522_t)
  );


  nor2s3
  U326
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n2523),
    .DIN2_t(n2523_t),
    .Q(WX9048),
    .Q_t(WX9048_t)
  );


  xor2s3
  U327
  (
    .DIN1(n5046),
    .DIN1_t(n5046_t),
    .DIN2(n3234),
    .DIN2_t(n3234_t),
    .Q(n2523),
    .Q_t(n2523_t)
  );


  nor2s3
  U328
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n2524),
    .DIN2_t(n2524_t),
    .Q(WX9046),
    .Q_t(WX9046_t)
  );


  xor2s3
  U329
  (
    .DIN1(n5042),
    .DIN1_t(n5042_t),
    .DIN2(n3233),
    .DIN2_t(n3233_t),
    .Q(n2524),
    .Q_t(n2524_t)
  );


  nor2s3
  U330
  (
    .DIN1(n2525),
    .DIN1_t(n2525_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX9044),
    .Q_t(WX9044_t)
  );


  xnr2s3
  U331
  (
    .DIN1(n3232),
    .DIN1_t(n3232_t),
    .DIN2(n2526),
    .DIN2_t(n2526_t),
    .Q(n2525),
    .Q_t(n2525_t)
  );


  xor2s3
  U332
  (
    .DIN1(n5038),
    .DIN1_t(n5038_t),
    .DIN2(n5122),
    .DIN2_t(n5122_t),
    .Q(n2526),
    .Q_t(n2526_t)
  );


  nor2s3
  U333
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n2527),
    .DIN2_t(n2527_t),
    .Q(WX9042),
    .Q_t(WX9042_t)
  );


  xor2s3
  U334
  (
    .DIN1(n5034),
    .DIN1_t(n5034_t),
    .DIN2(n3231),
    .DIN2_t(n3231_t),
    .Q(n2527),
    .Q_t(n2527_t)
  );


  nor2s3
  U335
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n2528),
    .DIN2_t(n2528_t),
    .Q(WX9040),
    .Q_t(WX9040_t)
  );


  xor2s3
  U336
  (
    .DIN1(n5030),
    .DIN1_t(n5030_t),
    .DIN2(n3230),
    .DIN2_t(n3230_t),
    .Q(n2528),
    .Q_t(n2528_t)
  );


  nor2s3
  U337
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n2529),
    .DIN2_t(n2529_t),
    .Q(WX9038),
    .Q_t(WX9038_t)
  );


  xor2s3
  U338
  (
    .DIN1(n5026),
    .DIN1_t(n5026_t),
    .DIN2(n3229),
    .DIN2_t(n3229_t),
    .Q(n2529),
    .Q_t(n2529_t)
  );


  nor2s3
  U339
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n2530),
    .DIN2_t(n2530_t),
    .Q(WX9036),
    .Q_t(WX9036_t)
  );


  xor2s3
  U340
  (
    .DIN1(n5022),
    .DIN1_t(n5022_t),
    .DIN2(n3228),
    .DIN2_t(n3228_t),
    .Q(n2530),
    .Q_t(n2530_t)
  );


  nor2s3
  U341
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n2531),
    .DIN2_t(n2531_t),
    .Q(WX9034),
    .Q_t(WX9034_t)
  );


  xor2s3
  U342
  (
    .DIN1(n5018),
    .DIN1_t(n5018_t),
    .DIN2(n3227),
    .DIN2_t(n3227_t),
    .Q(n2531),
    .Q_t(n2531_t)
  );


  nor2s3
  U343
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n2532),
    .DIN2_t(n2532_t),
    .Q(WX9032),
    .Q_t(WX9032_t)
  );


  xor2s3
  U344
  (
    .DIN1(n5014),
    .DIN1_t(n5014_t),
    .DIN2(n3226),
    .DIN2_t(n3226_t),
    .Q(n2532),
    .Q_t(n2532_t)
  );


  nor2s3
  U345
  (
    .DIN1(n2533),
    .DIN1_t(n2533_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX9030),
    .Q_t(WX9030_t)
  );


  xnr2s3
  U346
  (
    .DIN1(n3225),
    .DIN1_t(n3225_t),
    .DIN2(n2534),
    .DIN2_t(n2534_t),
    .Q(n2533),
    .Q_t(n2533_t)
  );


  xor2s3
  U347
  (
    .DIN1(n5010),
    .DIN1_t(n5010_t),
    .DIN2(n5122),
    .DIN2_t(n5122_t),
    .Q(n2534),
    .Q_t(n2534_t)
  );


  nor2s3
  U348
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n2535),
    .DIN2_t(n2535_t),
    .Q(WX9028),
    .Q_t(WX9028_t)
  );


  xor2s3
  U349
  (
    .DIN1(n5006),
    .DIN1_t(n5006_t),
    .DIN2(n3224),
    .DIN2_t(n3224_t),
    .Q(n2535),
    .Q_t(n2535_t)
  );


  nor2s3
  U350
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n2536),
    .DIN2_t(n2536_t),
    .Q(WX9026),
    .Q_t(WX9026_t)
  );


  xor2s3
  U351
  (
    .DIN1(n5002),
    .DIN1_t(n5002_t),
    .DIN2(n3223),
    .DIN2_t(n3223_t),
    .Q(n2536),
    .Q_t(n2536_t)
  );


  nor2s3
  U352
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n2537),
    .DIN2_t(n2537_t),
    .Q(WX9024),
    .Q_t(WX9024_t)
  );


  xor2s3
  U353
  (
    .DIN1(n4998),
    .DIN1_t(n4998_t),
    .DIN2(n3222),
    .DIN2_t(n3222_t),
    .Q(n2537),
    .Q_t(n2537_t)
  );


  nor2s3
  U354
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n2538),
    .DIN2_t(n2538_t),
    .Q(WX9022),
    .Q_t(WX9022_t)
  );


  xor2s3
  U355
  (
    .DIN1(n5122),
    .DIN1_t(n5122_t),
    .DIN2(n3221),
    .DIN2_t(n3221_t),
    .Q(n2538),
    .Q_t(n2538_t)
  );


  nor2s3
  U356
  (
    .DIN1(n6463),
    .DIN1_t(n6463_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX898),
    .Q_t(WX898_t)
  );


  nor2s3
  U357
  (
    .DIN1(n6527),
    .DIN1_t(n6527_t),
    .DIN2(n6737),
    .DIN2_t(n6737_t),
    .Q(WX896),
    .Q_t(WX896_t)
  );


  nor2s3
  U358
  (
    .DIN1(n6436),
    .DIN1_t(n6436_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX894),
    .Q_t(WX894_t)
  );


  nor2s3
  U359
  (
    .DIN1(n6469),
    .DIN1_t(n6469_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX892),
    .Q_t(WX892_t)
  );


  nor2s3
  U360
  (
    .DIN1(n6472),
    .DIN1_t(n6472_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX890),
    .Q_t(WX890_t)
  );


  nor2s3
  U361
  (
    .DIN1(n6460),
    .DIN1_t(n6460_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX888),
    .Q_t(WX888_t)
  );


  nor2s3
  U362
  (
    .DIN1(n6442),
    .DIN1_t(n6442_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX886),
    .Q_t(WX886_t)
  );


  nor2s3
  U363
  (
    .DIN1(n6466),
    .DIN1_t(n6466_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX884),
    .Q_t(WX884_t)
  );


  nor2s3
  U364
  (
    .DIN1(n6454),
    .DIN1_t(n6454_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX882),
    .Q_t(WX882_t)
  );


  nor2s3
  U365
  (
    .DIN1(n6504),
    .DIN1_t(n6504_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX880),
    .Q_t(WX880_t)
  );


  nor2s3
  U366
  (
    .DIN1(n6451),
    .DIN1_t(n6451_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX878),
    .Q_t(WX878_t)
  );


  nor2s3
  U367
  (
    .DIN1(n6445),
    .DIN1_t(n6445_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX876),
    .Q_t(WX876_t)
  );


  nor2s3
  U368
  (
    .DIN1(n6457),
    .DIN1_t(n6457_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX874),
    .Q_t(WX874_t)
  );


  nor2s3
  U369
  (
    .DIN1(n6448),
    .DIN1_t(n6448_t),
    .DIN2(n6736),
    .DIN2_t(n6736_t),
    .Q(WX872),
    .Q_t(WX872_t)
  );


  nor2s3
  U370
  (
    .DIN1(n6523),
    .DIN1_t(n6523_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX870),
    .Q_t(WX870_t)
  );


  nor2s3
  U371
  (
    .DIN1(n6439),
    .DIN1_t(n6439_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX868),
    .Q_t(WX868_t)
  );


  nor2s3
  U372
  (
    .DIN1(n6539),
    .DIN1_t(n6539_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX866),
    .Q_t(WX866_t)
  );


  nor2s3
  U373
  (
    .DIN1(n5157),
    .DIN1_t(n5157_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX8656),
    .Q_t(WX8656_t)
  );


  nor2s3
  U374
  (
    .DIN1(n5161),
    .DIN1_t(n5161_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX8654),
    .Q_t(WX8654_t)
  );


  nor2s3
  U375
  (
    .DIN1(n5165),
    .DIN1_t(n5165_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX8652),
    .Q_t(WX8652_t)
  );


  nor2s3
  U376
  (
    .DIN1(n5169),
    .DIN1_t(n5169_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX8650),
    .Q_t(WX8650_t)
  );


  nor2s3
  U377
  (
    .DIN1(n5173),
    .DIN1_t(n5173_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX8648),
    .Q_t(WX8648_t)
  );


  nor2s3
  U378
  (
    .DIN1(n5177),
    .DIN1_t(n5177_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX8646),
    .Q_t(WX8646_t)
  );


  nor2s3
  U379
  (
    .DIN1(n5181),
    .DIN1_t(n5181_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX8644),
    .Q_t(WX8644_t)
  );


  nor2s3
  U380
  (
    .DIN1(n5185),
    .DIN1_t(n5185_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX8642),
    .Q_t(WX8642_t)
  );


  nor2s3
  U381
  (
    .DIN1(n5189),
    .DIN1_t(n5189_t),
    .DIN2(n6735),
    .DIN2_t(n6735_t),
    .Q(WX8640),
    .Q_t(WX8640_t)
  );


  nor2s3
  U382
  (
    .DIN1(n6496),
    .DIN1_t(n6496_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX864),
    .Q_t(WX864_t)
  );


  nor2s3
  U383
  (
    .DIN1(n5193),
    .DIN1_t(n5193_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX8638),
    .Q_t(WX8638_t)
  );


  nor2s3
  U384
  (
    .DIN1(n5197),
    .DIN1_t(n5197_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX8636),
    .Q_t(WX8636_t)
  );


  nor2s3
  U385
  (
    .DIN1(n5201),
    .DIN1_t(n5201_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX8634),
    .Q_t(WX8634_t)
  );


  nor2s3
  U386
  (
    .DIN1(n5205),
    .DIN1_t(n5205_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX8632),
    .Q_t(WX8632_t)
  );


  nor2s3
  U387
  (
    .DIN1(n5209),
    .DIN1_t(n5209_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX8630),
    .Q_t(WX8630_t)
  );


  nor2s3
  U388
  (
    .DIN1(n5213),
    .DIN1_t(n5213_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX8628),
    .Q_t(WX8628_t)
  );


  nor2s3
  U389
  (
    .DIN1(n5217),
    .DIN1_t(n5217_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX8626),
    .Q_t(WX8626_t)
  );


  nor2s3
  U390
  (
    .DIN1(n5221),
    .DIN1_t(n5221_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX8624),
    .Q_t(WX8624_t)
  );


  nor2s3
  U391
  (
    .DIN1(n5226),
    .DIN1_t(n5226_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX8622),
    .Q_t(WX8622_t)
  );


  nor2s3
  U392
  (
    .DIN1(n5231),
    .DIN1_t(n5231_t),
    .DIN2(n6739),
    .DIN2_t(n6739_t),
    .Q(WX8620),
    .Q_t(WX8620_t)
  );


  nor2s3
  U393
  (
    .DIN1(n6544),
    .DIN1_t(n6544_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX862),
    .Q_t(WX862_t)
  );


  nor2s3
  U394
  (
    .DIN1(n5236),
    .DIN1_t(n5236_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX8618),
    .Q_t(WX8618_t)
  );


  nor2s3
  U395
  (
    .DIN1(n5241),
    .DIN1_t(n5241_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX8616),
    .Q_t(WX8616_t)
  );


  nor2s3
  U396
  (
    .DIN1(n5246),
    .DIN1_t(n5246_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX8614),
    .Q_t(WX8614_t)
  );


  nor2s3
  U397
  (
    .DIN1(n5251),
    .DIN1_t(n5251_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX8612),
    .Q_t(WX8612_t)
  );


  nor2s3
  U398
  (
    .DIN1(n5256),
    .DIN1_t(n5256_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX8610),
    .Q_t(WX8610_t)
  );


  nor2s3
  U399
  (
    .DIN1(n5261),
    .DIN1_t(n5261_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX8608),
    .Q_t(WX8608_t)
  );


  nor2s3
  U400
  (
    .DIN1(n5266),
    .DIN1_t(n5266_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX8606),
    .Q_t(WX8606_t)
  );


  nor2s3
  U401
  (
    .DIN1(n5271),
    .DIN1_t(n5271_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX8604),
    .Q_t(WX8604_t)
  );


  nor2s3
  U402
  (
    .DIN1(n5276),
    .DIN1_t(n5276_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX8602),
    .Q_t(WX8602_t)
  );


  nor2s3
  U403
  (
    .DIN1(n5281),
    .DIN1_t(n5281_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX8600),
    .Q_t(WX8600_t)
  );


  nor2s3
  U404
  (
    .DIN1(n6478),
    .DIN1_t(n6478_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX860),
    .Q_t(WX860_t)
  );


  nor2s3
  U405
  (
    .DIN1(n5286),
    .DIN1_t(n5286_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX8598),
    .Q_t(WX8598_t)
  );


  nor2s3
  U406
  (
    .DIN1(n5291),
    .DIN1_t(n5291_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX8596),
    .Q_t(WX8596_t)
  );


  nor2s3
  U407
  (
    .DIN1(n5296),
    .DIN1_t(n5296_t),
    .DIN2(n6755),
    .DIN2_t(n6755_t),
    .Q(WX8594),
    .Q_t(WX8594_t)
  );


  nor2s3
  U408
  (
    .DIN1(n5156),
    .DIN1_t(n5156_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX8592),
    .Q_t(WX8592_t)
  );


  nor2s3
  U409
  (
    .DIN1(n5160),
    .DIN1_t(n5160_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX8590),
    .Q_t(WX8590_t)
  );


  nor2s3
  U410
  (
    .DIN1(n5164),
    .DIN1_t(n5164_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX8588),
    .Q_t(WX8588_t)
  );


  nor2s3
  U411
  (
    .DIN1(n5168),
    .DIN1_t(n5168_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX8586),
    .Q_t(WX8586_t)
  );


  nor2s3
  U412
  (
    .DIN1(n5172),
    .DIN1_t(n5172_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX8584),
    .Q_t(WX8584_t)
  );


  nor2s3
  U413
  (
    .DIN1(n5176),
    .DIN1_t(n5176_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX8582),
    .Q_t(WX8582_t)
  );


  nor2s3
  U414
  (
    .DIN1(n5180),
    .DIN1_t(n5180_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX8580),
    .Q_t(WX8580_t)
  );


  nor2s3
  U415
  (
    .DIN1(n6535),
    .DIN1_t(n6535_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX858),
    .Q_t(WX858_t)
  );


  nor2s3
  U416
  (
    .DIN1(n5184),
    .DIN1_t(n5184_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX8578),
    .Q_t(WX8578_t)
  );


  nor2s3
  U417
  (
    .DIN1(n5188),
    .DIN1_t(n5188_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX8576),
    .Q_t(WX8576_t)
  );


  nor2s3
  U418
  (
    .DIN1(n5192),
    .DIN1_t(n5192_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX8574),
    .Q_t(WX8574_t)
  );


  nor2s3
  U419
  (
    .DIN1(n5196),
    .DIN1_t(n5196_t),
    .DIN2(n6754),
    .DIN2_t(n6754_t),
    .Q(WX8572),
    .Q_t(WX8572_t)
  );


  nor2s3
  U420
  (
    .DIN1(n5200),
    .DIN1_t(n5200_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX8570),
    .Q_t(WX8570_t)
  );


  nor2s3
  U421
  (
    .DIN1(n5204),
    .DIN1_t(n5204_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX8568),
    .Q_t(WX8568_t)
  );


  nor2s3
  U422
  (
    .DIN1(n5208),
    .DIN1_t(n5208_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX8566),
    .Q_t(WX8566_t)
  );


  nor2s3
  U423
  (
    .DIN1(n5212),
    .DIN1_t(n5212_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX8564),
    .Q_t(WX8564_t)
  );


  nor2s3
  U424
  (
    .DIN1(n5216),
    .DIN1_t(n5216_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX8562),
    .Q_t(WX8562_t)
  );


  and2s3
  U425
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5220),
    .DIN2_t(n5220_t),
    .Q(WX8560),
    .Q_t(WX8560_t)
  );


  nor2s3
  U426
  (
    .DIN1(n6518),
    .DIN1_t(n6518_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX856),
    .Q_t(WX856_t)
  );


  and2s3
  U427
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5225),
    .DIN2_t(n5225_t),
    .Q(WX8558),
    .Q_t(WX8558_t)
  );


  and2s3
  U428
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5230),
    .DIN2_t(n5230_t),
    .Q(WX8556),
    .Q_t(WX8556_t)
  );


  and2s3
  U429
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5235),
    .DIN2_t(n5235_t),
    .Q(WX8554),
    .Q_t(WX8554_t)
  );


  and2s3
  U430
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5240),
    .DIN2_t(n5240_t),
    .Q(WX8552),
    .Q_t(WX8552_t)
  );


  and2s3
  U431
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5245),
    .DIN2_t(n5245_t),
    .Q(WX8550),
    .Q_t(WX8550_t)
  );


  and2s3
  U432
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5250),
    .DIN2_t(n5250_t),
    .Q(WX8548),
    .Q_t(WX8548_t)
  );


  and2s3
  U433
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5255),
    .DIN2_t(n5255_t),
    .Q(WX8546),
    .Q_t(WX8546_t)
  );


  and2s3
  U434
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5260),
    .DIN2_t(n5260_t),
    .Q(WX8544),
    .Q_t(WX8544_t)
  );


  and2s3
  U435
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5265),
    .DIN2_t(n5265_t),
    .Q(WX8542),
    .Q_t(WX8542_t)
  );


  and2s3
  U436
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5270),
    .DIN2_t(n5270_t),
    .Q(WX8540),
    .Q_t(WX8540_t)
  );


  nor2s3
  U437
  (
    .DIN1(n6537),
    .DIN1_t(n6537_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX854),
    .Q_t(WX854_t)
  );


  and2s3
  U438
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5275),
    .DIN2_t(n5275_t),
    .Q(WX8538),
    .Q_t(WX8538_t)
  );


  and2s3
  U439
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5280),
    .DIN2_t(n5280_t),
    .Q(WX8536),
    .Q_t(WX8536_t)
  );


  and2s3
  U440
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5285),
    .DIN2_t(n5285_t),
    .Q(WX8534),
    .Q_t(WX8534_t)
  );


  and2s3
  U441
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5290),
    .DIN2_t(n5290_t),
    .Q(WX8532),
    .Q_t(WX8532_t)
  );


  and2s3
  U442
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5295),
    .DIN2_t(n5295_t),
    .Q(WX8530),
    .Q_t(WX8530_t)
  );


  and2s3
  U443
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5155),
    .DIN2_t(n5155_t),
    .Q(WX8528),
    .Q_t(WX8528_t)
  );


  and2s3
  U444
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5159),
    .DIN2_t(n5159_t),
    .Q(WX8526),
    .Q_t(WX8526_t)
  );


  and2s3
  U445
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5163),
    .DIN2_t(n5163_t),
    .Q(WX8524),
    .Q_t(WX8524_t)
  );


  and2s3
  U446
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5167),
    .DIN2_t(n5167_t),
    .Q(WX8522),
    .Q_t(WX8522_t)
  );


  and2s3
  U447
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5171),
    .DIN2_t(n5171_t),
    .Q(WX8520),
    .Q_t(WX8520_t)
  );


  nor2s3
  U448
  (
    .DIN1(n6512),
    .DIN1_t(n6512_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX852),
    .Q_t(WX852_t)
  );


  and2s3
  U449
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5175),
    .DIN2_t(n5175_t),
    .Q(WX8518),
    .Q_t(WX8518_t)
  );


  and2s3
  U450
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5179),
    .DIN2_t(n5179_t),
    .Q(WX8516),
    .Q_t(WX8516_t)
  );


  and2s3
  U451
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5183),
    .DIN2_t(n5183_t),
    .Q(WX8514),
    .Q_t(WX8514_t)
  );


  and2s3
  U452
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5187),
    .DIN2_t(n5187_t),
    .Q(WX8512),
    .Q_t(WX8512_t)
  );


  and2s3
  U453
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5191),
    .DIN2_t(n5191_t),
    .Q(WX8510),
    .Q_t(WX8510_t)
  );


  and2s3
  U454
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5195),
    .DIN2_t(n5195_t),
    .Q(WX8508),
    .Q_t(WX8508_t)
  );


  and2s3
  U455
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5199),
    .DIN2_t(n5199_t),
    .Q(WX8506),
    .Q_t(WX8506_t)
  );


  and2s3
  U456
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5203),
    .DIN2_t(n5203_t),
    .Q(WX8504),
    .Q_t(WX8504_t)
  );


  and2s3
  U457
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5207),
    .DIN2_t(n5207_t),
    .Q(WX8502),
    .Q_t(WX8502_t)
  );


  and2s3
  U458
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5211),
    .DIN2_t(n5211_t),
    .Q(WX8500),
    .Q_t(WX8500_t)
  );


  nor2s3
  U459
  (
    .DIN1(n6502),
    .DIN1_t(n6502_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX850),
    .Q_t(WX850_t)
  );


  and2s3
  U460
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5215),
    .DIN2_t(n5215_t),
    .Q(WX8498),
    .Q_t(WX8498_t)
  );


  nor2s3
  U461
  (
    .DIN1(n5219),
    .DIN1_t(n5219_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX8496),
    .Q_t(WX8496_t)
  );


  nor2s3
  U462
  (
    .DIN1(n5224),
    .DIN1_t(n5224_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX8494),
    .Q_t(WX8494_t)
  );


  nor2s3
  U463
  (
    .DIN1(n5229),
    .DIN1_t(n5229_t),
    .DIN2(n6753),
    .DIN2_t(n6753_t),
    .Q(WX8492),
    .Q_t(WX8492_t)
  );


  nor2s3
  U464
  (
    .DIN1(n5234),
    .DIN1_t(n5234_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX8490),
    .Q_t(WX8490_t)
  );


  nor2s3
  U465
  (
    .DIN1(n5239),
    .DIN1_t(n5239_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX8488),
    .Q_t(WX8488_t)
  );


  nor2s3
  U466
  (
    .DIN1(n5244),
    .DIN1_t(n5244_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX8486),
    .Q_t(WX8486_t)
  );


  nor2s3
  U467
  (
    .DIN1(n5249),
    .DIN1_t(n5249_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX8484),
    .Q_t(WX8484_t)
  );


  nor2s3
  U468
  (
    .DIN1(n5254),
    .DIN1_t(n5254_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX8482),
    .Q_t(WX8482_t)
  );


  nor2s3
  U469
  (
    .DIN1(n5259),
    .DIN1_t(n5259_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX8480),
    .Q_t(WX8480_t)
  );


  nor2s3
  U470
  (
    .DIN1(n6541),
    .DIN1_t(n6541_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX848),
    .Q_t(WX848_t)
  );


  nor2s3
  U471
  (
    .DIN1(n5264),
    .DIN1_t(n5264_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX8478),
    .Q_t(WX8478_t)
  );


  nor2s3
  U472
  (
    .DIN1(n5269),
    .DIN1_t(n5269_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX8476),
    .Q_t(WX8476_t)
  );


  nor2s3
  U473
  (
    .DIN1(n5274),
    .DIN1_t(n5274_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX8474),
    .Q_t(WX8474_t)
  );


  nor2s3
  U474
  (
    .DIN1(n5279),
    .DIN1_t(n5279_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX8472),
    .Q_t(WX8472_t)
  );


  nor2s3
  U475
  (
    .DIN1(n5284),
    .DIN1_t(n5284_t),
    .DIN2(n6752),
    .DIN2_t(n6752_t),
    .Q(WX8470),
    .Q_t(WX8470_t)
  );


  nor2s3
  U476
  (
    .DIN1(n5289),
    .DIN1_t(n5289_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX8468),
    .Q_t(WX8468_t)
  );


  nor2s3
  U477
  (
    .DIN1(n5294),
    .DIN1_t(n5294_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX8466),
    .Q_t(WX8466_t)
  );


  nnd4s2
  U478
  (
    .DIN1(n2539),
    .DIN1_t(n2539_t),
    .DIN2(n2540),
    .DIN2_t(n2540_t),
    .DIN3(n2541),
    .DIN3_t(n2541_t),
    .DIN4(n2542),
    .DIN4_t(n2542_t),
    .Q(WX8464),
    .Q_t(WX8464_t)
  );


  nnd2s3
  U479
  (
    .DIN1(n6625),
    .DIN1_t(n6625_t),
    .DIN2(n2313),
    .DIN2_t(n2313_t),
    .Q(n2542),
    .Q_t(n2542_t)
  );


  xor2s3
  U480
  (
    .DIN1(n2543),
    .DIN1_t(n2543_t),
    .DIN2(n2544),
    .DIN2_t(n2544_t),
    .Q(n2313),
    .Q_t(n2313_t)
  );


  xor2s3
  U481
  (
    .DIN1(n4995),
    .DIN1_t(n4995_t),
    .DIN2(n4996),
    .DIN2_t(n4996_t),
    .Q(n2544),
    .Q_t(n2544_t)
  );


  xnr2s3
  U482
  (
    .DIN1(n3205),
    .DIN1_t(n3205_t),
    .DIN2(n4997),
    .DIN2_t(n4997_t),
    .Q(n2543),
    .Q_t(n2543_t)
  );


  nnd2s3
  U483
  (
    .DIN1(n2545),
    .DIN1_t(n2545_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2541),
    .Q_t(n2541_t)
  );


  nnd2s3
  U484
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1889),
    .DIN2_t(n1889_t),
    .Q(n2540),
    .Q_t(n2540_t)
  );


  nnd2s3
  U485
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1888),
    .DIN2_t(n1888_t),
    .Q(n2539),
    .Q_t(n2539_t)
  );


  nnd4s2
  U486
  (
    .DIN1(n2546),
    .DIN1_t(n2546_t),
    .DIN2(n2547),
    .DIN2_t(n2547_t),
    .DIN3(n2548),
    .DIN3_t(n2548_t),
    .DIN4(n2549),
    .DIN4_t(n2549_t),
    .Q(WX8462),
    .Q_t(WX8462_t)
  );


  nnd2s3
  U487
  (
    .DIN1(n2322),
    .DIN1_t(n2322_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2549),
    .Q_t(n2549_t)
  );


  xor2s3
  U488
  (
    .DIN1(n2550),
    .DIN1_t(n2550_t),
    .DIN2(n2551),
    .DIN2_t(n2551_t),
    .Q(n2322),
    .Q_t(n2322_t)
  );


  xor2s3
  U489
  (
    .DIN1(n4999),
    .DIN1_t(n4999_t),
    .DIN2(n5000),
    .DIN2_t(n5000_t),
    .Q(n2551),
    .Q_t(n2551_t)
  );


  xnr2s3
  U490
  (
    .DIN1(n3206),
    .DIN1_t(n3206_t),
    .DIN2(n5001),
    .DIN2_t(n5001_t),
    .Q(n2550),
    .Q_t(n2550_t)
  );


  nnd2s3
  U491
  (
    .DIN1(n2552),
    .DIN1_t(n2552_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2548),
    .Q_t(n2548_t)
  );


  nnd2s3
  U492
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1890),
    .DIN2_t(n1890_t),
    .Q(n2547),
    .Q_t(n2547_t)
  );


  nnd2s3
  U493
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1887),
    .DIN2_t(n1887_t),
    .Q(n2546),
    .Q_t(n2546_t)
  );


  nnd4s2
  U494
  (
    .DIN1(n2553),
    .DIN1_t(n2553_t),
    .DIN2(n2554),
    .DIN2_t(n2554_t),
    .DIN3(n2555),
    .DIN3_t(n2555_t),
    .DIN4(n2556),
    .DIN4_t(n2556_t),
    .Q(WX8460),
    .Q_t(WX8460_t)
  );


  nnd2s3
  U495
  (
    .DIN1(n2328),
    .DIN1_t(n2328_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2556),
    .Q_t(n2556_t)
  );


  xor2s3
  U496
  (
    .DIN1(n2557),
    .DIN1_t(n2557_t),
    .DIN2(n2558),
    .DIN2_t(n2558_t),
    .Q(n2328),
    .Q_t(n2328_t)
  );


  xor2s3
  U497
  (
    .DIN1(n5003),
    .DIN1_t(n5003_t),
    .DIN2(n5004),
    .DIN2_t(n5004_t),
    .Q(n2558),
    .Q_t(n2558_t)
  );


  xnr2s3
  U498
  (
    .DIN1(n3207),
    .DIN1_t(n3207_t),
    .DIN2(n5005),
    .DIN2_t(n5005_t),
    .Q(n2557),
    .Q_t(n2557_t)
  );


  nnd2s3
  U499
  (
    .DIN1(n2559),
    .DIN1_t(n2559_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2555),
    .Q_t(n2555_t)
  );


  nnd2s3
  U500
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1891),
    .DIN2_t(n1891_t),
    .Q(n2554),
    .Q_t(n2554_t)
  );


  nnd2s3
  U501
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1886),
    .DIN2_t(n1886_t),
    .Q(n2553),
    .Q_t(n2553_t)
  );


  nor2s3
  U502
  (
    .DIN1(n6493),
    .DIN1_t(n6493_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX846),
    .Q_t(WX846_t)
  );


  nnd4s2
  U503
  (
    .DIN1(n2560),
    .DIN1_t(n2560_t),
    .DIN2(n2561),
    .DIN2_t(n2561_t),
    .DIN3(n2562),
    .DIN3_t(n2562_t),
    .DIN4(n2563),
    .DIN4_t(n2563_t),
    .Q(WX8458),
    .Q_t(WX8458_t)
  );


  nnd2s3
  U504
  (
    .DIN1(n2334),
    .DIN1_t(n2334_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2563),
    .Q_t(n2563_t)
  );


  xor2s3
  U505
  (
    .DIN1(n2564),
    .DIN1_t(n2564_t),
    .DIN2(n2565),
    .DIN2_t(n2565_t),
    .Q(n2334),
    .Q_t(n2334_t)
  );


  xor2s3
  U506
  (
    .DIN1(n5007),
    .DIN1_t(n5007_t),
    .DIN2(n5008),
    .DIN2_t(n5008_t),
    .Q(n2565),
    .Q_t(n2565_t)
  );


  xnr2s3
  U507
  (
    .DIN1(n3208),
    .DIN1_t(n3208_t),
    .DIN2(n5009),
    .DIN2_t(n5009_t),
    .Q(n2564),
    .Q_t(n2564_t)
  );


  nnd2s3
  U508
  (
    .DIN1(n2566),
    .DIN1_t(n2566_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2562),
    .Q_t(n2562_t)
  );


  nnd2s3
  U509
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1892),
    .DIN2_t(n1892_t),
    .Q(n2561),
    .Q_t(n2561_t)
  );


  nnd2s3
  U510
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1885),
    .DIN2_t(n1885_t),
    .Q(n2560),
    .Q_t(n2560_t)
  );


  nnd4s2
  U511
  (
    .DIN1(n2567),
    .DIN1_t(n2567_t),
    .DIN2(n2568),
    .DIN2_t(n2568_t),
    .DIN3(n2569),
    .DIN3_t(n2569_t),
    .DIN4(n2570),
    .DIN4_t(n2570_t),
    .Q(WX8456),
    .Q_t(WX8456_t)
  );


  nnd2s3
  U512
  (
    .DIN1(n2340),
    .DIN1_t(n2340_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2570),
    .Q_t(n2570_t)
  );


  xor2s3
  U513
  (
    .DIN1(n2571),
    .DIN1_t(n2571_t),
    .DIN2(n2572),
    .DIN2_t(n2572_t),
    .Q(n2340),
    .Q_t(n2340_t)
  );


  xor2s3
  U514
  (
    .DIN1(n5011),
    .DIN1_t(n5011_t),
    .DIN2(n5012),
    .DIN2_t(n5012_t),
    .Q(n2572),
    .Q_t(n2572_t)
  );


  xnr2s3
  U515
  (
    .DIN1(n3209),
    .DIN1_t(n3209_t),
    .DIN2(n5013),
    .DIN2_t(n5013_t),
    .Q(n2571),
    .Q_t(n2571_t)
  );


  nnd2s3
  U516
  (
    .DIN1(n2573),
    .DIN1_t(n2573_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2569),
    .Q_t(n2569_t)
  );


  nnd2s3
  U517
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1893),
    .DIN2_t(n1893_t),
    .Q(n2568),
    .Q_t(n2568_t)
  );


  nnd2s3
  U518
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1884),
    .DIN2_t(n1884_t),
    .Q(n2567),
    .Q_t(n2567_t)
  );


  nnd4s2
  U519
  (
    .DIN1(n2574),
    .DIN1_t(n2574_t),
    .DIN2(n2575),
    .DIN2_t(n2575_t),
    .DIN3(n2576),
    .DIN3_t(n2576_t),
    .DIN4(n2577),
    .DIN4_t(n2577_t),
    .Q(WX8454),
    .Q_t(WX8454_t)
  );


  nnd2s3
  U520
  (
    .DIN1(n2346),
    .DIN1_t(n2346_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2577),
    .Q_t(n2577_t)
  );


  xor2s3
  U521
  (
    .DIN1(n2578),
    .DIN1_t(n2578_t),
    .DIN2(n2579),
    .DIN2_t(n2579_t),
    .Q(n2346),
    .Q_t(n2346_t)
  );


  xor2s3
  U522
  (
    .DIN1(n5015),
    .DIN1_t(n5015_t),
    .DIN2(n5016),
    .DIN2_t(n5016_t),
    .Q(n2579),
    .Q_t(n2579_t)
  );


  xnr2s3
  U523
  (
    .DIN1(n3210),
    .DIN1_t(n3210_t),
    .DIN2(n5017),
    .DIN2_t(n5017_t),
    .Q(n2578),
    .Q_t(n2578_t)
  );


  nnd2s3
  U524
  (
    .DIN1(n2580),
    .DIN1_t(n2580_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2576),
    .Q_t(n2576_t)
  );


  nnd2s3
  U525
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1894),
    .DIN2_t(n1894_t),
    .Q(n2575),
    .Q_t(n2575_t)
  );


  nnd2s3
  U526
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1883),
    .DIN2_t(n1883_t),
    .Q(n2574),
    .Q_t(n2574_t)
  );


  nnd4s2
  U527
  (
    .DIN1(n2581),
    .DIN1_t(n2581_t),
    .DIN2(n2582),
    .DIN2_t(n2582_t),
    .DIN3(n2583),
    .DIN3_t(n2583_t),
    .DIN4(n2584),
    .DIN4_t(n2584_t),
    .Q(WX8452),
    .Q_t(WX8452_t)
  );


  nnd2s3
  U528
  (
    .DIN1(n2352),
    .DIN1_t(n2352_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2584),
    .Q_t(n2584_t)
  );


  xor2s3
  U529
  (
    .DIN1(n2585),
    .DIN1_t(n2585_t),
    .DIN2(n2586),
    .DIN2_t(n2586_t),
    .Q(n2352),
    .Q_t(n2352_t)
  );


  xor2s3
  U530
  (
    .DIN1(n5019),
    .DIN1_t(n5019_t),
    .DIN2(n5020),
    .DIN2_t(n5020_t),
    .Q(n2586),
    .Q_t(n2586_t)
  );


  xnr2s3
  U531
  (
    .DIN1(n3211),
    .DIN1_t(n3211_t),
    .DIN2(n5021),
    .DIN2_t(n5021_t),
    .Q(n2585),
    .Q_t(n2585_t)
  );


  nnd2s3
  U532
  (
    .DIN1(n2587),
    .DIN1_t(n2587_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2583),
    .Q_t(n2583_t)
  );


  nnd2s3
  U533
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1895),
    .DIN2_t(n1895_t),
    .Q(n2582),
    .Q_t(n2582_t)
  );


  nnd2s3
  U534
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1882),
    .DIN2_t(n1882_t),
    .Q(n2581),
    .Q_t(n2581_t)
  );


  nnd4s2
  U535
  (
    .DIN1(n2588),
    .DIN1_t(n2588_t),
    .DIN2(n2589),
    .DIN2_t(n2589_t),
    .DIN3(n2590),
    .DIN3_t(n2590_t),
    .DIN4(n2591),
    .DIN4_t(n2591_t),
    .Q(WX8450),
    .Q_t(WX8450_t)
  );


  nnd2s3
  U536
  (
    .DIN1(n2358),
    .DIN1_t(n2358_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2591),
    .Q_t(n2591_t)
  );


  xor2s3
  U537
  (
    .DIN1(n2592),
    .DIN1_t(n2592_t),
    .DIN2(n2593),
    .DIN2_t(n2593_t),
    .Q(n2358),
    .Q_t(n2358_t)
  );


  xor2s3
  U538
  (
    .DIN1(n5023),
    .DIN1_t(n5023_t),
    .DIN2(n5024),
    .DIN2_t(n5024_t),
    .Q(n2593),
    .Q_t(n2593_t)
  );


  xnr2s3
  U539
  (
    .DIN1(n3212),
    .DIN1_t(n3212_t),
    .DIN2(n5025),
    .DIN2_t(n5025_t),
    .Q(n2592),
    .Q_t(n2592_t)
  );


  nnd2s3
  U540
  (
    .DIN1(n2594),
    .DIN1_t(n2594_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2590),
    .Q_t(n2590_t)
  );


  nnd2s3
  U541
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1896),
    .DIN2_t(n1896_t),
    .Q(n2589),
    .Q_t(n2589_t)
  );


  nnd2s3
  U542
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1881),
    .DIN2_t(n1881_t),
    .Q(n2588),
    .Q_t(n2588_t)
  );


  nnd4s2
  U543
  (
    .DIN1(n2595),
    .DIN1_t(n2595_t),
    .DIN2(n2596),
    .DIN2_t(n2596_t),
    .DIN3(n2597),
    .DIN3_t(n2597_t),
    .DIN4(n2598),
    .DIN4_t(n2598_t),
    .Q(WX8448),
    .Q_t(WX8448_t)
  );


  nnd2s3
  U544
  (
    .DIN1(n2364),
    .DIN1_t(n2364_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2598),
    .Q_t(n2598_t)
  );


  xor2s3
  U545
  (
    .DIN1(n2599),
    .DIN1_t(n2599_t),
    .DIN2(n2600),
    .DIN2_t(n2600_t),
    .Q(n2364),
    .Q_t(n2364_t)
  );


  xor2s3
  U546
  (
    .DIN1(n5027),
    .DIN1_t(n5027_t),
    .DIN2(n5028),
    .DIN2_t(n5028_t),
    .Q(n2600),
    .Q_t(n2600_t)
  );


  xnr2s3
  U547
  (
    .DIN1(n3213),
    .DIN1_t(n3213_t),
    .DIN2(n5029),
    .DIN2_t(n5029_t),
    .Q(n2599),
    .Q_t(n2599_t)
  );


  nnd2s3
  U548
  (
    .DIN1(n2601),
    .DIN1_t(n2601_t),
    .DIN2(n6664),
    .DIN2_t(n6664_t),
    .Q(n2597),
    .Q_t(n2597_t)
  );


  nnd2s3
  U549
  (
    .DIN1(n6613),
    .DIN1_t(n6613_t),
    .DIN2(n1897),
    .DIN2_t(n1897_t),
    .Q(n2596),
    .Q_t(n2596_t)
  );


  nnd2s3
  U550
  (
    .DIN1(n6582),
    .DIN1_t(n6582_t),
    .DIN2(n1880),
    .DIN2_t(n1880_t),
    .Q(n2595),
    .Q_t(n2595_t)
  );


  nnd4s2
  U551
  (
    .DIN1(n2602),
    .DIN1_t(n2602_t),
    .DIN2(n2603),
    .DIN2_t(n2603_t),
    .DIN3(n2604),
    .DIN3_t(n2604_t),
    .DIN4(n2605),
    .DIN4_t(n2605_t),
    .Q(WX8446),
    .Q_t(WX8446_t)
  );


  nnd2s3
  U552
  (
    .DIN1(n2370),
    .DIN1_t(n2370_t),
    .DIN2(n6633),
    .DIN2_t(n6633_t),
    .Q(n2605),
    .Q_t(n2605_t)
  );


  xor2s3
  U553
  (
    .DIN1(n2606),
    .DIN1_t(n2606_t),
    .DIN2(n2607),
    .DIN2_t(n2607_t),
    .Q(n2370),
    .Q_t(n2370_t)
  );


  xor2s3
  U554
  (
    .DIN1(n5031),
    .DIN1_t(n5031_t),
    .DIN2(n5032),
    .DIN2_t(n5032_t),
    .Q(n2607),
    .Q_t(n2607_t)
  );


  xnr2s3
  U555
  (
    .DIN1(n3214),
    .DIN1_t(n3214_t),
    .DIN2(n5033),
    .DIN2_t(n5033_t),
    .Q(n2606),
    .Q_t(n2606_t)
  );


  nnd2s3
  U556
  (
    .DIN1(n2608),
    .DIN1_t(n2608_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2604),
    .Q_t(n2604_t)
  );


  nnd2s3
  U557
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1898),
    .DIN2_t(n1898_t),
    .Q(n2603),
    .Q_t(n2603_t)
  );


  nnd2s3
  U558
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1879),
    .DIN2_t(n1879_t),
    .Q(n2602),
    .Q_t(n2602_t)
  );


  nnd4s2
  U559
  (
    .DIN1(n2609),
    .DIN1_t(n2609_t),
    .DIN2(n2610),
    .DIN2_t(n2610_t),
    .DIN3(n2611),
    .DIN3_t(n2611_t),
    .DIN4(n2612),
    .DIN4_t(n2612_t),
    .Q(WX8444),
    .Q_t(WX8444_t)
  );


  nnd2s3
  U560
  (
    .DIN1(n2376),
    .DIN1_t(n2376_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2612),
    .Q_t(n2612_t)
  );


  xor2s3
  U561
  (
    .DIN1(n2613),
    .DIN1_t(n2613_t),
    .DIN2(n2614),
    .DIN2_t(n2614_t),
    .Q(n2376),
    .Q_t(n2376_t)
  );


  xor2s3
  U562
  (
    .DIN1(n5035),
    .DIN1_t(n5035_t),
    .DIN2(n5036),
    .DIN2_t(n5036_t),
    .Q(n2614),
    .Q_t(n2614_t)
  );


  xnr2s3
  U563
  (
    .DIN1(n3215),
    .DIN1_t(n3215_t),
    .DIN2(n5037),
    .DIN2_t(n5037_t),
    .Q(n2613),
    .Q_t(n2613_t)
  );


  nnd2s3
  U564
  (
    .DIN1(n2615),
    .DIN1_t(n2615_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2611),
    .Q_t(n2611_t)
  );


  nnd2s3
  U565
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1899),
    .DIN2_t(n1899_t),
    .Q(n2610),
    .Q_t(n2610_t)
  );


  nnd2s3
  U566
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1878),
    .DIN2_t(n1878_t),
    .Q(n2609),
    .Q_t(n2609_t)
  );


  nnd4s2
  U567
  (
    .DIN1(n2616),
    .DIN1_t(n2616_t),
    .DIN2(n2617),
    .DIN2_t(n2617_t),
    .DIN3(n2618),
    .DIN3_t(n2618_t),
    .DIN4(n2619),
    .DIN4_t(n2619_t),
    .Q(WX8442),
    .Q_t(WX8442_t)
  );


  nnd2s3
  U568
  (
    .DIN1(n2382),
    .DIN1_t(n2382_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2619),
    .Q_t(n2619_t)
  );


  xor2s3
  U569
  (
    .DIN1(n2620),
    .DIN1_t(n2620_t),
    .DIN2(n2621),
    .DIN2_t(n2621_t),
    .Q(n2382),
    .Q_t(n2382_t)
  );


  xor2s3
  U570
  (
    .DIN1(n5039),
    .DIN1_t(n5039_t),
    .DIN2(n5040),
    .DIN2_t(n5040_t),
    .Q(n2621),
    .Q_t(n2621_t)
  );


  xnr2s3
  U571
  (
    .DIN1(n3216),
    .DIN1_t(n3216_t),
    .DIN2(n5041),
    .DIN2_t(n5041_t),
    .Q(n2620),
    .Q_t(n2620_t)
  );


  nnd2s3
  U572
  (
    .DIN1(n2622),
    .DIN1_t(n2622_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2618),
    .Q_t(n2618_t)
  );


  nnd2s3
  U573
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1900),
    .DIN2_t(n1900_t),
    .Q(n2617),
    .Q_t(n2617_t)
  );


  nnd2s3
  U574
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1877),
    .DIN2_t(n1877_t),
    .Q(n2616),
    .Q_t(n2616_t)
  );


  nnd4s2
  U575
  (
    .DIN1(n2623),
    .DIN1_t(n2623_t),
    .DIN2(n2624),
    .DIN2_t(n2624_t),
    .DIN3(n2625),
    .DIN3_t(n2625_t),
    .DIN4(n2626),
    .DIN4_t(n2626_t),
    .Q(WX8440),
    .Q_t(WX8440_t)
  );


  nnd2s3
  U576
  (
    .DIN1(n2388),
    .DIN1_t(n2388_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2626),
    .Q_t(n2626_t)
  );


  xor2s3
  U577
  (
    .DIN1(n2627),
    .DIN1_t(n2627_t),
    .DIN2(n2628),
    .DIN2_t(n2628_t),
    .Q(n2388),
    .Q_t(n2388_t)
  );


  xor2s3
  U578
  (
    .DIN1(n5043),
    .DIN1_t(n5043_t),
    .DIN2(n5044),
    .DIN2_t(n5044_t),
    .Q(n2628),
    .Q_t(n2628_t)
  );


  xnr2s3
  U579
  (
    .DIN1(n3217),
    .DIN1_t(n3217_t),
    .DIN2(n5045),
    .DIN2_t(n5045_t),
    .Q(n2627),
    .Q_t(n2627_t)
  );


  nnd2s3
  U580
  (
    .DIN1(n2629),
    .DIN1_t(n2629_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2625),
    .Q_t(n2625_t)
  );


  nnd2s3
  U581
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1901),
    .DIN2_t(n1901_t),
    .Q(n2624),
    .Q_t(n2624_t)
  );


  nnd2s3
  U582
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1876),
    .DIN2_t(n1876_t),
    .Q(n2623),
    .Q_t(n2623_t)
  );


  nor2s3
  U583
  (
    .DIN1(n6487),
    .DIN1_t(n6487_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX844),
    .Q_t(WX844_t)
  );


  nnd4s2
  U584
  (
    .DIN1(n2630),
    .DIN1_t(n2630_t),
    .DIN2(n2631),
    .DIN2_t(n2631_t),
    .DIN3(n2632),
    .DIN3_t(n2632_t),
    .DIN4(n2633),
    .DIN4_t(n2633_t),
    .Q(WX8438),
    .Q_t(WX8438_t)
  );


  nnd2s3
  U585
  (
    .DIN1(n2394),
    .DIN1_t(n2394_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2633),
    .Q_t(n2633_t)
  );


  xor2s3
  U586
  (
    .DIN1(n2634),
    .DIN1_t(n2634_t),
    .DIN2(n2635),
    .DIN2_t(n2635_t),
    .Q(n2394),
    .Q_t(n2394_t)
  );


  xor2s3
  U587
  (
    .DIN1(n5047),
    .DIN1_t(n5047_t),
    .DIN2(n5048),
    .DIN2_t(n5048_t),
    .Q(n2635),
    .Q_t(n2635_t)
  );


  xnr2s3
  U588
  (
    .DIN1(n3218),
    .DIN1_t(n3218_t),
    .DIN2(n5049),
    .DIN2_t(n5049_t),
    .Q(n2634),
    .Q_t(n2634_t)
  );


  nnd2s3
  U589
  (
    .DIN1(n2636),
    .DIN1_t(n2636_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2632),
    .Q_t(n2632_t)
  );


  nnd2s3
  U590
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1902),
    .DIN2_t(n1902_t),
    .Q(n2631),
    .Q_t(n2631_t)
  );


  nnd2s3
  U591
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1875),
    .DIN2_t(n1875_t),
    .Q(n2630),
    .Q_t(n2630_t)
  );


  nnd4s2
  U592
  (
    .DIN1(n2637),
    .DIN1_t(n2637_t),
    .DIN2(n2638),
    .DIN2_t(n2638_t),
    .DIN3(n2639),
    .DIN3_t(n2639_t),
    .DIN4(n2640),
    .DIN4_t(n2640_t),
    .Q(WX8436),
    .Q_t(WX8436_t)
  );


  nnd2s3
  U593
  (
    .DIN1(n2400),
    .DIN1_t(n2400_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2640),
    .Q_t(n2640_t)
  );


  xor2s3
  U594
  (
    .DIN1(n2641),
    .DIN1_t(n2641_t),
    .DIN2(n2642),
    .DIN2_t(n2642_t),
    .Q(n2400),
    .Q_t(n2400_t)
  );


  xor2s3
  U595
  (
    .DIN1(n5051),
    .DIN1_t(n5051_t),
    .DIN2(n5052),
    .DIN2_t(n5052_t),
    .Q(n2642),
    .Q_t(n2642_t)
  );


  xnr2s3
  U596
  (
    .DIN1(n3219),
    .DIN1_t(n3219_t),
    .DIN2(n5053),
    .DIN2_t(n5053_t),
    .Q(n2641),
    .Q_t(n2641_t)
  );


  nnd2s3
  U597
  (
    .DIN1(n2643),
    .DIN1_t(n2643_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2639),
    .Q_t(n2639_t)
  );


  nnd2s3
  U598
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1903),
    .DIN2_t(n1903_t),
    .Q(n2638),
    .Q_t(n2638_t)
  );


  nnd2s3
  U599
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1874),
    .DIN2_t(n1874_t),
    .Q(n2637),
    .Q_t(n2637_t)
  );


  nnd4s2
  U600
  (
    .DIN1(n2644),
    .DIN1_t(n2644_t),
    .DIN2(n2645),
    .DIN2_t(n2645_t),
    .DIN3(n2646),
    .DIN3_t(n2646_t),
    .DIN4(n2647),
    .DIN4_t(n2647_t),
    .Q(WX8434),
    .Q_t(WX8434_t)
  );


  nnd2s3
  U601
  (
    .DIN1(n2406),
    .DIN1_t(n2406_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2647),
    .Q_t(n2647_t)
  );


  xor2s3
  U602
  (
    .DIN1(n2648),
    .DIN1_t(n2648_t),
    .DIN2(n2649),
    .DIN2_t(n2649_t),
    .Q(n2406),
    .Q_t(n2406_t)
  );


  xor2s3
  U603
  (
    .DIN1(n5055),
    .DIN1_t(n5055_t),
    .DIN2(n5056),
    .DIN2_t(n5056_t),
    .Q(n2649),
    .Q_t(n2649_t)
  );


  xnr2s3
  U604
  (
    .DIN1(n3220),
    .DIN1_t(n3220_t),
    .DIN2(n5057),
    .DIN2_t(n5057_t),
    .Q(n2648),
    .Q_t(n2648_t)
  );


  nnd2s3
  U605
  (
    .DIN1(n2650),
    .DIN1_t(n2650_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2646),
    .Q_t(n2646_t)
  );


  nnd2s3
  U606
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1904),
    .DIN2_t(n1904_t),
    .Q(n2645),
    .Q_t(n2645_t)
  );


  nnd2s3
  U607
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1873),
    .DIN2_t(n1873_t),
    .Q(n2644),
    .Q_t(n2644_t)
  );


  nnd4s2
  U608
  (
    .DIN1(n2651),
    .DIN1_t(n2651_t),
    .DIN2(n2652),
    .DIN2_t(n2652_t),
    .DIN3(n2653),
    .DIN3_t(n2653_t),
    .DIN4(n2654),
    .DIN4_t(n2654_t),
    .Q(WX8432),
    .Q_t(WX8432_t)
  );


  nnd2s3
  U609
  (
    .DIN1(n2412),
    .DIN1_t(n2412_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2654),
    .Q_t(n2654_t)
  );


  xor2s3
  U610
  (
    .DIN1(n2655),
    .DIN1_t(n2655_t),
    .DIN2(n2656),
    .DIN2_t(n2656_t),
    .Q(n2412),
    .Q_t(n2412_t)
  );


  xor2s3
  U611
  (
    .DIN1(n5061),
    .DIN1_t(n5061_t),
    .DIN2(n2657),
    .DIN2_t(n2657_t),
    .Q(n2656),
    .Q_t(n2656_t)
  );


  xor2s3
  U612
  (
    .DIN1(n5059),
    .DIN1_t(n5059_t),
    .DIN2(n5060),
    .DIN2_t(n5060_t),
    .Q(n2657),
    .Q_t(n2657_t)
  );


  xor2s3
  U613
  (
    .DIN1(n6414),
    .DIN1_t(n6414_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n2655),
    .Q_t(n2655_t)
  );


  nnd2s3
  U614
  (
    .DIN1(n2658),
    .DIN1_t(n2658_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2653),
    .Q_t(n2653_t)
  );


  nnd2s3
  U615
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1905),
    .DIN2_t(n1905_t),
    .Q(n2652),
    .Q_t(n2652_t)
  );


  nnd2s3
  U616
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1872),
    .DIN2_t(n1872_t),
    .Q(n2651),
    .Q_t(n2651_t)
  );


  nnd4s2
  U617
  (
    .DIN1(n2659),
    .DIN1_t(n2659_t),
    .DIN2(n2660),
    .DIN2_t(n2660_t),
    .DIN3(n2661),
    .DIN3_t(n2661_t),
    .DIN4(n2662),
    .DIN4_t(n2662_t),
    .Q(WX8430),
    .Q_t(WX8430_t)
  );


  nnd2s3
  U618
  (
    .DIN1(n2418),
    .DIN1_t(n2418_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2662),
    .Q_t(n2662_t)
  );


  xor2s3
  U619
  (
    .DIN1(n2663),
    .DIN1_t(n2663_t),
    .DIN2(n2664),
    .DIN2_t(n2664_t),
    .Q(n2418),
    .Q_t(n2418_t)
  );


  xor2s3
  U620
  (
    .DIN1(n5065),
    .DIN1_t(n5065_t),
    .DIN2(n2665),
    .DIN2_t(n2665_t),
    .Q(n2664),
    .Q_t(n2664_t)
  );


  xor2s3
  U621
  (
    .DIN1(n5063),
    .DIN1_t(n5063_t),
    .DIN2(n5064),
    .DIN2_t(n5064_t),
    .Q(n2665),
    .Q_t(n2665_t)
  );


  xor2s3
  U622
  (
    .DIN1(n6412),
    .DIN1_t(n6412_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2663),
    .Q_t(n2663_t)
  );


  nnd2s3
  U623
  (
    .DIN1(n2666),
    .DIN1_t(n2666_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2661),
    .Q_t(n2661_t)
  );


  nnd2s3
  U624
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1906),
    .DIN2_t(n1906_t),
    .Q(n2660),
    .Q_t(n2660_t)
  );


  nnd2s3
  U625
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1871),
    .DIN2_t(n1871_t),
    .Q(n2659),
    .Q_t(n2659_t)
  );


  nnd4s2
  U626
  (
    .DIN1(n2667),
    .DIN1_t(n2667_t),
    .DIN2(n2668),
    .DIN2_t(n2668_t),
    .DIN3(n2669),
    .DIN3_t(n2669_t),
    .DIN4(n2670),
    .DIN4_t(n2670_t),
    .Q(WX8428),
    .Q_t(WX8428_t)
  );


  nnd2s3
  U627
  (
    .DIN1(n2424),
    .DIN1_t(n2424_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2670),
    .Q_t(n2670_t)
  );


  xor2s3
  U628
  (
    .DIN1(n2671),
    .DIN1_t(n2671_t),
    .DIN2(n2672),
    .DIN2_t(n2672_t),
    .Q(n2424),
    .Q_t(n2424_t)
  );


  xor2s3
  U629
  (
    .DIN1(n5069),
    .DIN1_t(n5069_t),
    .DIN2(n2673),
    .DIN2_t(n2673_t),
    .Q(n2672),
    .Q_t(n2672_t)
  );


  xor2s3
  U630
  (
    .DIN1(n5067),
    .DIN1_t(n5067_t),
    .DIN2(n5068),
    .DIN2_t(n5068_t),
    .Q(n2673),
    .Q_t(n2673_t)
  );


  xor2s3
  U631
  (
    .DIN1(n6410),
    .DIN1_t(n6410_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2671),
    .Q_t(n2671_t)
  );


  nnd2s3
  U632
  (
    .DIN1(n2674),
    .DIN1_t(n2674_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2669),
    .Q_t(n2669_t)
  );


  nnd2s3
  U633
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1907),
    .DIN2_t(n1907_t),
    .Q(n2668),
    .Q_t(n2668_t)
  );


  nnd2s3
  U634
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1870),
    .DIN2_t(n1870_t),
    .Q(n2667),
    .Q_t(n2667_t)
  );


  nnd4s2
  U635
  (
    .DIN1(n2675),
    .DIN1_t(n2675_t),
    .DIN2(n2676),
    .DIN2_t(n2676_t),
    .DIN3(n2677),
    .DIN3_t(n2677_t),
    .DIN4(n2678),
    .DIN4_t(n2678_t),
    .Q(WX8426),
    .Q_t(WX8426_t)
  );


  nnd2s3
  U636
  (
    .DIN1(n2430),
    .DIN1_t(n2430_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2678),
    .Q_t(n2678_t)
  );


  xor2s3
  U637
  (
    .DIN1(n2679),
    .DIN1_t(n2679_t),
    .DIN2(n2680),
    .DIN2_t(n2680_t),
    .Q(n2430),
    .Q_t(n2430_t)
  );


  xor2s3
  U638
  (
    .DIN1(n5073),
    .DIN1_t(n5073_t),
    .DIN2(n2681),
    .DIN2_t(n2681_t),
    .Q(n2680),
    .Q_t(n2680_t)
  );


  xor2s3
  U639
  (
    .DIN1(n5071),
    .DIN1_t(n5071_t),
    .DIN2(n5072),
    .DIN2_t(n5072_t),
    .Q(n2681),
    .Q_t(n2681_t)
  );


  xor2s3
  U640
  (
    .DIN1(n6408),
    .DIN1_t(n6408_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2679),
    .Q_t(n2679_t)
  );


  nnd2s3
  U641
  (
    .DIN1(n2682),
    .DIN1_t(n2682_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2677),
    .Q_t(n2677_t)
  );


  nnd2s3
  U642
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1908),
    .DIN2_t(n1908_t),
    .Q(n2676),
    .Q_t(n2676_t)
  );


  nnd2s3
  U643
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1869),
    .DIN2_t(n1869_t),
    .Q(n2675),
    .Q_t(n2675_t)
  );


  nnd4s2
  U644
  (
    .DIN1(n2683),
    .DIN1_t(n2683_t),
    .DIN2(n2684),
    .DIN2_t(n2684_t),
    .DIN3(n2685),
    .DIN3_t(n2685_t),
    .DIN4(n2686),
    .DIN4_t(n2686_t),
    .Q(WX8424),
    .Q_t(WX8424_t)
  );


  nnd2s3
  U645
  (
    .DIN1(n2436),
    .DIN1_t(n2436_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2686),
    .Q_t(n2686_t)
  );


  xor2s3
  U646
  (
    .DIN1(n2687),
    .DIN1_t(n2687_t),
    .DIN2(n2688),
    .DIN2_t(n2688_t),
    .Q(n2436),
    .Q_t(n2436_t)
  );


  xor2s3
  U647
  (
    .DIN1(n5077),
    .DIN1_t(n5077_t),
    .DIN2(n2689),
    .DIN2_t(n2689_t),
    .Q(n2688),
    .Q_t(n2688_t)
  );


  xor2s3
  U648
  (
    .DIN1(n5075),
    .DIN1_t(n5075_t),
    .DIN2(n5076),
    .DIN2_t(n5076_t),
    .Q(n2689),
    .Q_t(n2689_t)
  );


  xor2s3
  U649
  (
    .DIN1(n6406),
    .DIN1_t(n6406_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2687),
    .Q_t(n2687_t)
  );


  nnd2s3
  U650
  (
    .DIN1(n2690),
    .DIN1_t(n2690_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2685),
    .Q_t(n2685_t)
  );


  nnd2s3
  U651
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1909),
    .DIN2_t(n1909_t),
    .Q(n2684),
    .Q_t(n2684_t)
  );


  nnd2s3
  U652
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1868),
    .DIN2_t(n1868_t),
    .Q(n2683),
    .Q_t(n2683_t)
  );


  nnd4s2
  U653
  (
    .DIN1(n2691),
    .DIN1_t(n2691_t),
    .DIN2(n2692),
    .DIN2_t(n2692_t),
    .DIN3(n2693),
    .DIN3_t(n2693_t),
    .DIN4(n2694),
    .DIN4_t(n2694_t),
    .Q(WX8422),
    .Q_t(WX8422_t)
  );


  nnd2s3
  U654
  (
    .DIN1(n2442),
    .DIN1_t(n2442_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2694),
    .Q_t(n2694_t)
  );


  xor2s3
  U655
  (
    .DIN1(n2695),
    .DIN1_t(n2695_t),
    .DIN2(n2696),
    .DIN2_t(n2696_t),
    .Q(n2442),
    .Q_t(n2442_t)
  );


  xor2s3
  U656
  (
    .DIN1(n5081),
    .DIN1_t(n5081_t),
    .DIN2(n2697),
    .DIN2_t(n2697_t),
    .Q(n2696),
    .Q_t(n2696_t)
  );


  xor2s3
  U657
  (
    .DIN1(n5079),
    .DIN1_t(n5079_t),
    .DIN2(n5080),
    .DIN2_t(n5080_t),
    .Q(n2697),
    .Q_t(n2697_t)
  );


  xor2s3
  U658
  (
    .DIN1(n6404),
    .DIN1_t(n6404_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2695),
    .Q_t(n2695_t)
  );


  nnd2s3
  U659
  (
    .DIN1(n2698),
    .DIN1_t(n2698_t),
    .DIN2(n6663),
    .DIN2_t(n6663_t),
    .Q(n2693),
    .Q_t(n2693_t)
  );


  nnd2s3
  U660
  (
    .DIN1(n6612),
    .DIN1_t(n6612_t),
    .DIN2(n1910),
    .DIN2_t(n1910_t),
    .Q(n2692),
    .Q_t(n2692_t)
  );


  nnd2s3
  U661
  (
    .DIN1(n6581),
    .DIN1_t(n6581_t),
    .DIN2(n1867),
    .DIN2_t(n1867_t),
    .Q(n2691),
    .Q_t(n2691_t)
  );


  nnd4s2
  U662
  (
    .DIN1(n2699),
    .DIN1_t(n2699_t),
    .DIN2(n2700),
    .DIN2_t(n2700_t),
    .DIN3(n2701),
    .DIN3_t(n2701_t),
    .DIN4(n2702),
    .DIN4_t(n2702_t),
    .Q(WX8420),
    .Q_t(WX8420_t)
  );


  nnd2s3
  U663
  (
    .DIN1(n2448),
    .DIN1_t(n2448_t),
    .DIN2(n6632),
    .DIN2_t(n6632_t),
    .Q(n2702),
    .Q_t(n2702_t)
  );


  xor2s3
  U664
  (
    .DIN1(n2703),
    .DIN1_t(n2703_t),
    .DIN2(n2704),
    .DIN2_t(n2704_t),
    .Q(n2448),
    .Q_t(n2448_t)
  );


  xor2s3
  U665
  (
    .DIN1(n5085),
    .DIN1_t(n5085_t),
    .DIN2(n2705),
    .DIN2_t(n2705_t),
    .Q(n2704),
    .Q_t(n2704_t)
  );


  xor2s3
  U666
  (
    .DIN1(n5083),
    .DIN1_t(n5083_t),
    .DIN2(n5084),
    .DIN2_t(n5084_t),
    .Q(n2705),
    .Q_t(n2705_t)
  );


  xor2s3
  U667
  (
    .DIN1(n6402),
    .DIN1_t(n6402_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2703),
    .Q_t(n2703_t)
  );


  nnd2s3
  U668
  (
    .DIN1(n2706),
    .DIN1_t(n2706_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2701),
    .Q_t(n2701_t)
  );


  nnd2s3
  U669
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1911),
    .DIN2_t(n1911_t),
    .Q(n2700),
    .Q_t(n2700_t)
  );


  nnd2s3
  U670
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1866),
    .DIN2_t(n1866_t),
    .Q(n2699),
    .Q_t(n2699_t)
  );


  nor2s3
  U671
  (
    .DIN1(n6484),
    .DIN1_t(n6484_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX842),
    .Q_t(WX842_t)
  );


  nnd4s2
  U672
  (
    .DIN1(n2707),
    .DIN1_t(n2707_t),
    .DIN2(n2708),
    .DIN2_t(n2708_t),
    .DIN3(n2709),
    .DIN3_t(n2709_t),
    .DIN4(n2710),
    .DIN4_t(n2710_t),
    .Q(WX8418),
    .Q_t(WX8418_t)
  );


  nnd2s3
  U673
  (
    .DIN1(n2454),
    .DIN1_t(n2454_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2710),
    .Q_t(n2710_t)
  );


  xor2s3
  U674
  (
    .DIN1(n2711),
    .DIN1_t(n2711_t),
    .DIN2(n2712),
    .DIN2_t(n2712_t),
    .Q(n2454),
    .Q_t(n2454_t)
  );


  xor2s3
  U675
  (
    .DIN1(n5089),
    .DIN1_t(n5089_t),
    .DIN2(n2713),
    .DIN2_t(n2713_t),
    .Q(n2712),
    .Q_t(n2712_t)
  );


  xor2s3
  U676
  (
    .DIN1(n5087),
    .DIN1_t(n5087_t),
    .DIN2(n5088),
    .DIN2_t(n5088_t),
    .Q(n2713),
    .Q_t(n2713_t)
  );


  xor2s3
  U677
  (
    .DIN1(n6400),
    .DIN1_t(n6400_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2711),
    .Q_t(n2711_t)
  );


  nnd2s3
  U678
  (
    .DIN1(n2714),
    .DIN1_t(n2714_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2709),
    .Q_t(n2709_t)
  );


  nnd2s3
  U679
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1912),
    .DIN2_t(n1912_t),
    .Q(n2708),
    .Q_t(n2708_t)
  );


  nnd2s3
  U680
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1865),
    .DIN2_t(n1865_t),
    .Q(n2707),
    .Q_t(n2707_t)
  );


  nnd4s2
  U681
  (
    .DIN1(n2715),
    .DIN1_t(n2715_t),
    .DIN2(n2716),
    .DIN2_t(n2716_t),
    .DIN3(n2717),
    .DIN3_t(n2717_t),
    .DIN4(n2718),
    .DIN4_t(n2718_t),
    .Q(WX8416),
    .Q_t(WX8416_t)
  );


  nnd2s3
  U682
  (
    .DIN1(n2460),
    .DIN1_t(n2460_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2718),
    .Q_t(n2718_t)
  );


  xor2s3
  U683
  (
    .DIN1(n2719),
    .DIN1_t(n2719_t),
    .DIN2(n2720),
    .DIN2_t(n2720_t),
    .Q(n2460),
    .Q_t(n2460_t)
  );


  xor2s3
  U684
  (
    .DIN1(n5093),
    .DIN1_t(n5093_t),
    .DIN2(n2721),
    .DIN2_t(n2721_t),
    .Q(n2720),
    .Q_t(n2720_t)
  );


  xor2s3
  U685
  (
    .DIN1(n5091),
    .DIN1_t(n5091_t),
    .DIN2(n5092),
    .DIN2_t(n5092_t),
    .Q(n2721),
    .Q_t(n2721_t)
  );


  xor2s3
  U686
  (
    .DIN1(n6398),
    .DIN1_t(n6398_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2719),
    .Q_t(n2719_t)
  );


  nnd2s3
  U687
  (
    .DIN1(n2722),
    .DIN1_t(n2722_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2717),
    .Q_t(n2717_t)
  );


  nnd2s3
  U688
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1913),
    .DIN2_t(n1913_t),
    .Q(n2716),
    .Q_t(n2716_t)
  );


  nnd2s3
  U689
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1864),
    .DIN2_t(n1864_t),
    .Q(n2715),
    .Q_t(n2715_t)
  );


  nnd4s2
  U690
  (
    .DIN1(n2723),
    .DIN1_t(n2723_t),
    .DIN2(n2724),
    .DIN2_t(n2724_t),
    .DIN3(n2725),
    .DIN3_t(n2725_t),
    .DIN4(n2726),
    .DIN4_t(n2726_t),
    .Q(WX8414),
    .Q_t(WX8414_t)
  );


  nnd2s3
  U691
  (
    .DIN1(n2466),
    .DIN1_t(n2466_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2726),
    .Q_t(n2726_t)
  );


  xor2s3
  U692
  (
    .DIN1(n2727),
    .DIN1_t(n2727_t),
    .DIN2(n2728),
    .DIN2_t(n2728_t),
    .Q(n2466),
    .Q_t(n2466_t)
  );


  xor2s3
  U693
  (
    .DIN1(n5097),
    .DIN1_t(n5097_t),
    .DIN2(n2729),
    .DIN2_t(n2729_t),
    .Q(n2728),
    .Q_t(n2728_t)
  );


  xor2s3
  U694
  (
    .DIN1(n5095),
    .DIN1_t(n5095_t),
    .DIN2(n5096),
    .DIN2_t(n5096_t),
    .Q(n2729),
    .Q_t(n2729_t)
  );


  xor2s3
  U695
  (
    .DIN1(n6396),
    .DIN1_t(n6396_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2727),
    .Q_t(n2727_t)
  );


  nnd2s3
  U696
  (
    .DIN1(n2730),
    .DIN1_t(n2730_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2725),
    .Q_t(n2725_t)
  );


  nnd2s3
  U697
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1914),
    .DIN2_t(n1914_t),
    .Q(n2724),
    .Q_t(n2724_t)
  );


  nnd2s3
  U698
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1863),
    .DIN2_t(n1863_t),
    .Q(n2723),
    .Q_t(n2723_t)
  );


  nnd4s2
  U699
  (
    .DIN1(n2731),
    .DIN1_t(n2731_t),
    .DIN2(n2732),
    .DIN2_t(n2732_t),
    .DIN3(n2733),
    .DIN3_t(n2733_t),
    .DIN4(n2734),
    .DIN4_t(n2734_t),
    .Q(WX8412),
    .Q_t(WX8412_t)
  );


  nnd2s3
  U700
  (
    .DIN1(n2472),
    .DIN1_t(n2472_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2734),
    .Q_t(n2734_t)
  );


  xor2s3
  U701
  (
    .DIN1(n2735),
    .DIN1_t(n2735_t),
    .DIN2(n2736),
    .DIN2_t(n2736_t),
    .Q(n2472),
    .Q_t(n2472_t)
  );


  xor2s3
  U702
  (
    .DIN1(n5101),
    .DIN1_t(n5101_t),
    .DIN2(n2737),
    .DIN2_t(n2737_t),
    .Q(n2736),
    .Q_t(n2736_t)
  );


  xor2s3
  U703
  (
    .DIN1(n5099),
    .DIN1_t(n5099_t),
    .DIN2(n5100),
    .DIN2_t(n5100_t),
    .Q(n2737),
    .Q_t(n2737_t)
  );


  xor2s3
  U704
  (
    .DIN1(n6394),
    .DIN1_t(n6394_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2735),
    .Q_t(n2735_t)
  );


  nnd2s3
  U705
  (
    .DIN1(n2738),
    .DIN1_t(n2738_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2733),
    .Q_t(n2733_t)
  );


  nnd2s3
  U706
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1915),
    .DIN2_t(n1915_t),
    .Q(n2732),
    .Q_t(n2732_t)
  );


  nnd2s3
  U707
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1862),
    .DIN2_t(n1862_t),
    .Q(n2731),
    .Q_t(n2731_t)
  );


  nnd4s2
  U708
  (
    .DIN1(n2739),
    .DIN1_t(n2739_t),
    .DIN2(n2740),
    .DIN2_t(n2740_t),
    .DIN3(n2741),
    .DIN3_t(n2741_t),
    .DIN4(n2742),
    .DIN4_t(n2742_t),
    .Q(WX8410),
    .Q_t(WX8410_t)
  );


  nnd2s3
  U709
  (
    .DIN1(n2478),
    .DIN1_t(n2478_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2742),
    .Q_t(n2742_t)
  );


  xor2s3
  U710
  (
    .DIN1(n2743),
    .DIN1_t(n2743_t),
    .DIN2(n2744),
    .DIN2_t(n2744_t),
    .Q(n2478),
    .Q_t(n2478_t)
  );


  xor2s3
  U711
  (
    .DIN1(n5105),
    .DIN1_t(n5105_t),
    .DIN2(n2745),
    .DIN2_t(n2745_t),
    .Q(n2744),
    .Q_t(n2744_t)
  );


  xor2s3
  U712
  (
    .DIN1(n5103),
    .DIN1_t(n5103_t),
    .DIN2(n5104),
    .DIN2_t(n5104_t),
    .Q(n2745),
    .Q_t(n2745_t)
  );


  xor2s3
  U713
  (
    .DIN1(n6392),
    .DIN1_t(n6392_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2743),
    .Q_t(n2743_t)
  );


  nnd2s3
  U714
  (
    .DIN1(n2746),
    .DIN1_t(n2746_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2741),
    .Q_t(n2741_t)
  );


  nnd2s3
  U715
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1916),
    .DIN2_t(n1916_t),
    .Q(n2740),
    .Q_t(n2740_t)
  );


  nnd2s3
  U716
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1861),
    .DIN2_t(n1861_t),
    .Q(n2739),
    .Q_t(n2739_t)
  );


  nnd4s2
  U717
  (
    .DIN1(n2747),
    .DIN1_t(n2747_t),
    .DIN2(n2748),
    .DIN2_t(n2748_t),
    .DIN3(n2749),
    .DIN3_t(n2749_t),
    .DIN4(n2750),
    .DIN4_t(n2750_t),
    .Q(WX8408),
    .Q_t(WX8408_t)
  );


  nnd2s3
  U718
  (
    .DIN1(n2484),
    .DIN1_t(n2484_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2750),
    .Q_t(n2750_t)
  );


  xor2s3
  U719
  (
    .DIN1(n2751),
    .DIN1_t(n2751_t),
    .DIN2(n2752),
    .DIN2_t(n2752_t),
    .Q(n2484),
    .Q_t(n2484_t)
  );


  xor2s3
  U720
  (
    .DIN1(n5109),
    .DIN1_t(n5109_t),
    .DIN2(n2753),
    .DIN2_t(n2753_t),
    .Q(n2752),
    .Q_t(n2752_t)
  );


  xor2s3
  U721
  (
    .DIN1(n5107),
    .DIN1_t(n5107_t),
    .DIN2(n5108),
    .DIN2_t(n5108_t),
    .Q(n2753),
    .Q_t(n2753_t)
  );


  xor2s3
  U722
  (
    .DIN1(n6390),
    .DIN1_t(n6390_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n2751),
    .Q_t(n2751_t)
  );


  nnd2s3
  U723
  (
    .DIN1(n2754),
    .DIN1_t(n2754_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2749),
    .Q_t(n2749_t)
  );


  nnd2s3
  U724
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1917),
    .DIN2_t(n1917_t),
    .Q(n2748),
    .Q_t(n2748_t)
  );


  nnd2s3
  U725
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1860),
    .DIN2_t(n1860_t),
    .Q(n2747),
    .Q_t(n2747_t)
  );


  nnd4s2
  U726
  (
    .DIN1(n2755),
    .DIN1_t(n2755_t),
    .DIN2(n2756),
    .DIN2_t(n2756_t),
    .DIN3(n2757),
    .DIN3_t(n2757_t),
    .DIN4(n2758),
    .DIN4_t(n2758_t),
    .Q(WX8406),
    .Q_t(WX8406_t)
  );


  nnd2s3
  U727
  (
    .DIN1(n2490),
    .DIN1_t(n2490_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2758),
    .Q_t(n2758_t)
  );


  xor2s3
  U728
  (
    .DIN1(n2759),
    .DIN1_t(n2759_t),
    .DIN2(n2760),
    .DIN2_t(n2760_t),
    .Q(n2490),
    .Q_t(n2490_t)
  );


  xor2s3
  U729
  (
    .DIN1(n5113),
    .DIN1_t(n5113_t),
    .DIN2(n2761),
    .DIN2_t(n2761_t),
    .Q(n2760),
    .Q_t(n2760_t)
  );


  xor2s3
  U730
  (
    .DIN1(n5111),
    .DIN1_t(n5111_t),
    .DIN2(n5112),
    .DIN2_t(n5112_t),
    .Q(n2761),
    .Q_t(n2761_t)
  );


  xor2s3
  U731
  (
    .DIN1(n6388),
    .DIN1_t(n6388_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2759),
    .Q_t(n2759_t)
  );


  nnd2s3
  U732
  (
    .DIN1(n2762),
    .DIN1_t(n2762_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2757),
    .Q_t(n2757_t)
  );


  nnd2s3
  U733
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1918),
    .DIN2_t(n1918_t),
    .Q(n2756),
    .Q_t(n2756_t)
  );


  nnd2s3
  U734
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1859),
    .DIN2_t(n1859_t),
    .Q(n2755),
    .Q_t(n2755_t)
  );


  nnd4s2
  U735
  (
    .DIN1(n2763),
    .DIN1_t(n2763_t),
    .DIN2(n2764),
    .DIN2_t(n2764_t),
    .DIN3(n2765),
    .DIN3_t(n2765_t),
    .DIN4(n2766),
    .DIN4_t(n2766_t),
    .Q(WX8404),
    .Q_t(WX8404_t)
  );


  nnd2s3
  U736
  (
    .DIN1(n2496),
    .DIN1_t(n2496_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2766),
    .Q_t(n2766_t)
  );


  xor2s3
  U737
  (
    .DIN1(n2767),
    .DIN1_t(n2767_t),
    .DIN2(n2768),
    .DIN2_t(n2768_t),
    .Q(n2496),
    .Q_t(n2496_t)
  );


  xor2s3
  U738
  (
    .DIN1(n5117),
    .DIN1_t(n5117_t),
    .DIN2(n2769),
    .DIN2_t(n2769_t),
    .Q(n2768),
    .Q_t(n2768_t)
  );


  xor2s3
  U739
  (
    .DIN1(n5115),
    .DIN1_t(n5115_t),
    .DIN2(n5116),
    .DIN2_t(n5116_t),
    .Q(n2769),
    .Q_t(n2769_t)
  );


  xor2s3
  U740
  (
    .DIN1(n6386),
    .DIN1_t(n6386_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2767),
    .Q_t(n2767_t)
  );


  nnd2s3
  U741
  (
    .DIN1(n2770),
    .DIN1_t(n2770_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2765),
    .Q_t(n2765_t)
  );


  nnd2s3
  U742
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1919),
    .DIN2_t(n1919_t),
    .Q(n2764),
    .Q_t(n2764_t)
  );


  nnd2s3
  U743
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1858),
    .DIN2_t(n1858_t),
    .Q(n2763),
    .Q_t(n2763_t)
  );


  nnd4s2
  U744
  (
    .DIN1(n2771),
    .DIN1_t(n2771_t),
    .DIN2(n2772),
    .DIN2_t(n2772_t),
    .DIN3(n2773),
    .DIN3_t(n2773_t),
    .DIN4(n2774),
    .DIN4_t(n2774_t),
    .Q(WX8402),
    .Q_t(WX8402_t)
  );


  nnd2s3
  U745
  (
    .DIN1(n2502),
    .DIN1_t(n2502_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2774),
    .Q_t(n2774_t)
  );


  xor2s3
  U746
  (
    .DIN1(n2775),
    .DIN1_t(n2775_t),
    .DIN2(n2776),
    .DIN2_t(n2776_t),
    .Q(n2502),
    .Q_t(n2502_t)
  );


  xor2s3
  U747
  (
    .DIN1(n5121),
    .DIN1_t(n5121_t),
    .DIN2(n2777),
    .DIN2_t(n2777_t),
    .Q(n2776),
    .Q_t(n2776_t)
  );


  xor2s3
  U748
  (
    .DIN1(n5119),
    .DIN1_t(n5119_t),
    .DIN2(n5120),
    .DIN2_t(n5120_t),
    .Q(n2777),
    .Q_t(n2777_t)
  );


  xor2s3
  U749
  (
    .DIN1(n6384),
    .DIN1_t(n6384_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2775),
    .Q_t(n2775_t)
  );


  nnd2s3
  U750
  (
    .DIN1(n2778),
    .DIN1_t(n2778_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2773),
    .Q_t(n2773_t)
  );


  nnd2s3
  U751
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1920),
    .DIN2_t(n1920_t),
    .Q(n2772),
    .Q_t(n2772_t)
  );


  nnd2s3
  U752
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1857),
    .DIN2_t(n1857_t),
    .Q(n2771),
    .Q_t(n2771_t)
  );


  nor2s3
  U753
  (
    .DIN1(n6547),
    .DIN1_t(n6547_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX840),
    .Q_t(WX840_t)
  );


  nor2s3
  U754
  (
    .DIN1(n6475),
    .DIN1_t(n6475_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX838),
    .Q_t(WX838_t)
  );


  nor2s3
  U755
  (
    .DIN1(n6531),
    .DIN1_t(n6531_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX836),
    .Q_t(WX836_t)
  );


  nor2s3
  U756
  (
    .DIN1(n6464),
    .DIN1_t(n6464_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX834),
    .Q_t(WX834_t)
  );


  nor2s3
  U757
  (
    .DIN1(n6528),
    .DIN1_t(n6528_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX832),
    .Q_t(WX832_t)
  );


  nor2s3
  U758
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n1920),
    .DIN2_t(n1920_t),
    .Q(WX8304),
    .Q_t(WX8304_t)
  );


  nor2s3
  U759
  (
    .DIN1(n5124),
    .DIN1_t(n5124_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX8302),
    .Q_t(WX8302_t)
  );


  nor2s3
  U760
  (
    .DIN1(n5125),
    .DIN1_t(n5125_t),
    .DIN2(n6751),
    .DIN2_t(n6751_t),
    .Q(WX8300),
    .Q_t(WX8300_t)
  );


  nor2s3
  U761
  (
    .DIN1(n6562),
    .DIN1_t(n6562_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX830),
    .Q_t(WX830_t)
  );


  nor2s3
  U762
  (
    .DIN1(n5126),
    .DIN1_t(n5126_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX8298),
    .Q_t(WX8298_t)
  );


  nor2s3
  U763
  (
    .DIN1(n5127),
    .DIN1_t(n5127_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX8296),
    .Q_t(WX8296_t)
  );


  nor2s3
  U764
  (
    .DIN1(n5128),
    .DIN1_t(n5128_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX8294),
    .Q_t(WX8294_t)
  );


  nor2s3
  U765
  (
    .DIN1(n5129),
    .DIN1_t(n5129_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX8292),
    .Q_t(WX8292_t)
  );


  nor2s3
  U766
  (
    .DIN1(n5130),
    .DIN1_t(n5130_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX8290),
    .Q_t(WX8290_t)
  );


  nor2s3
  U767
  (
    .DIN1(n5131),
    .DIN1_t(n5131_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX8288),
    .Q_t(WX8288_t)
  );


  nor2s3
  U768
  (
    .DIN1(n5132),
    .DIN1_t(n5132_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX8286),
    .Q_t(WX8286_t)
  );


  nor2s3
  U769
  (
    .DIN1(n5133),
    .DIN1_t(n5133_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX8284),
    .Q_t(WX8284_t)
  );


  nor2s3
  U770
  (
    .DIN1(n5134),
    .DIN1_t(n5134_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX8282),
    .Q_t(WX8282_t)
  );


  nor2s3
  U771
  (
    .DIN1(n5135),
    .DIN1_t(n5135_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX8280),
    .Q_t(WX8280_t)
  );


  nor2s3
  U772
  (
    .DIN1(n6470),
    .DIN1_t(n6470_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX828),
    .Q_t(WX828_t)
  );


  nor2s3
  U773
  (
    .DIN1(n5136),
    .DIN1_t(n5136_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX8278),
    .Q_t(WX8278_t)
  );


  nor2s3
  U774
  (
    .DIN1(n5137),
    .DIN1_t(n5137_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX8276),
    .Q_t(WX8276_t)
  );


  nor2s3
  U775
  (
    .DIN1(n5138),
    .DIN1_t(n5138_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX8274),
    .Q_t(WX8274_t)
  );


  nor2s3
  U776
  (
    .DIN1(n5139),
    .DIN1_t(n5139_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX8272),
    .Q_t(WX8272_t)
  );


  nor2s3
  U777
  (
    .DIN1(n5140),
    .DIN1_t(n5140_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX8270),
    .Q_t(WX8270_t)
  );


  nor2s3
  U778
  (
    .DIN1(n5141),
    .DIN1_t(n5141_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX8268),
    .Q_t(WX8268_t)
  );


  nor2s3
  U779
  (
    .DIN1(n5142),
    .DIN1_t(n5142_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX8266),
    .Q_t(WX8266_t)
  );


  nor2s3
  U780
  (
    .DIN1(n5143),
    .DIN1_t(n5143_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX8264),
    .Q_t(WX8264_t)
  );


  nor2s3
  U781
  (
    .DIN1(n5144),
    .DIN1_t(n5144_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX8262),
    .Q_t(WX8262_t)
  );


  nor2s3
  U782
  (
    .DIN1(n5145),
    .DIN1_t(n5145_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX8260),
    .Q_t(WX8260_t)
  );


  nor2s3
  U783
  (
    .DIN1(n6473),
    .DIN1_t(n6473_t),
    .DIN2(n6749),
    .DIN2_t(n6749_t),
    .Q(WX826),
    .Q_t(WX826_t)
  );


  nor2s3
  U784
  (
    .DIN1(n5146),
    .DIN1_t(n5146_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX8258),
    .Q_t(WX8258_t)
  );


  nor2s3
  U785
  (
    .DIN1(n5147),
    .DIN1_t(n5147_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX8256),
    .Q_t(WX8256_t)
  );


  nor2s3
  U786
  (
    .DIN1(n5148),
    .DIN1_t(n5148_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX8254),
    .Q_t(WX8254_t)
  );


  nor2s3
  U787
  (
    .DIN1(n5149),
    .DIN1_t(n5149_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX8252),
    .Q_t(WX8252_t)
  );


  nor2s3
  U788
  (
    .DIN1(n5150),
    .DIN1_t(n5150_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX8250),
    .Q_t(WX8250_t)
  );


  nor2s3
  U789
  (
    .DIN1(n5151),
    .DIN1_t(n5151_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX8248),
    .Q_t(WX8248_t)
  );


  nor2s3
  U790
  (
    .DIN1(n5152),
    .DIN1_t(n5152_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX8246),
    .Q_t(WX8246_t)
  );


  nor2s3
  U791
  (
    .DIN1(n5153),
    .DIN1_t(n5153_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX8244),
    .Q_t(WX8244_t)
  );


  nor2s3
  U792
  (
    .DIN1(n5154),
    .DIN1_t(n5154_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX8242),
    .Q_t(WX8242_t)
  );


  nor2s3
  U793
  (
    .DIN1(n6461),
    .DIN1_t(n6461_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX824),
    .Q_t(WX824_t)
  );


  nor2s3
  U794
  (
    .DIN1(n6443),
    .DIN1_t(n6443_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX822),
    .Q_t(WX822_t)
  );


  nor2s3
  U795
  (
    .DIN1(n6467),
    .DIN1_t(n6467_t),
    .DIN2(n6748),
    .DIN2_t(n6748_t),
    .Q(WX820),
    .Q_t(WX820_t)
  );


  nor2s3
  U796
  (
    .DIN1(n6455),
    .DIN1_t(n6455_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX818),
    .Q_t(WX818_t)
  );


  nor2s3
  U797
  (
    .DIN1(n6505),
    .DIN1_t(n6505_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX816),
    .Q_t(WX816_t)
  );


  nor2s3
  U798
  (
    .DIN1(n6452),
    .DIN1_t(n6452_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX814),
    .Q_t(WX814_t)
  );


  nor2s3
  U799
  (
    .DIN1(n6446),
    .DIN1_t(n6446_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX812),
    .Q_t(WX812_t)
  );


  nor2s3
  U800
  (
    .DIN1(n6458),
    .DIN1_t(n6458_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX810),
    .Q_t(WX810_t)
  );


  nor2s3
  U801
  (
    .DIN1(n6449),
    .DIN1_t(n6449_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX808),
    .Q_t(WX808_t)
  );


  nor2s3
  U802
  (
    .DIN1(n6524),
    .DIN1_t(n6524_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX806),
    .Q_t(WX806_t)
  );


  nor2s3
  U803
  (
    .DIN1(n6440),
    .DIN1_t(n6440_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX804),
    .Q_t(WX804_t)
  );


  nor2s3
  U804
  (
    .DIN1(n6508),
    .DIN1_t(n6508_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX802),
    .Q_t(WX802_t)
  );


  nor2s3
  U805
  (
    .DIN1(n6497),
    .DIN1_t(n6497_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX800),
    .Q_t(WX800_t)
  );


  nor2s3
  U806
  (
    .DIN1(n6489),
    .DIN1_t(n6489_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX798),
    .Q_t(WX798_t)
  );


  nor2s3
  U807
  (
    .DIN1(n6479),
    .DIN1_t(n6479_t),
    .DIN2(n6747),
    .DIN2_t(n6747_t),
    .Q(WX796),
    .Q_t(WX796_t)
  );


  nor2s3
  U808
  (
    .DIN1(n6520),
    .DIN1_t(n6520_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX794),
    .Q_t(WX794_t)
  );


  nor2s3
  U809
  (
    .DIN1(n6519),
    .DIN1_t(n6519_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX792),
    .Q_t(WX792_t)
  );


  nor2s3
  U810
  (
    .DIN1(n6514),
    .DIN1_t(n6514_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX790),
    .Q_t(WX790_t)
  );


  nor2s3
  U811
  (
    .DIN1(n6513),
    .DIN1_t(n6513_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX788),
    .Q_t(WX788_t)
  );


  nor2s3
  U812
  (
    .DIN1(n6503),
    .DIN1_t(n6503_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX786),
    .Q_t(WX786_t)
  );


  nor2s3
  U813
  (
    .DIN1(n6498),
    .DIN1_t(n6498_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX784),
    .Q_t(WX784_t)
  );


  nor2s3
  U814
  (
    .DIN1(n6494),
    .DIN1_t(n6494_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX782),
    .Q_t(WX782_t)
  );


  nor2s3
  U815
  (
    .DIN1(n6488),
    .DIN1_t(n6488_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX780),
    .Q_t(WX780_t)
  );


  nor2s3
  U816
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n2779),
    .DIN2_t(n2779_t),
    .Q(WX7791),
    .Q_t(WX7791_t)
  );


  xor2s3
  U817
  (
    .DIN1(n5293),
    .DIN1_t(n5293_t),
    .DIN2(n5473),
    .DIN2_t(n5473_t),
    .Q(n2779),
    .Q_t(n2779_t)
  );


  nor2s3
  U818
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n2780),
    .DIN2_t(n2780_t),
    .Q(WX7789),
    .Q_t(WX7789_t)
  );


  xor2s3
  U819
  (
    .DIN1(n5288),
    .DIN1_t(n5288_t),
    .DIN2(n5468),
    .DIN2_t(n5468_t),
    .Q(n2780),
    .Q_t(n2780_t)
  );


  nor2s3
  U820
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n2781),
    .DIN2_t(n2781_t),
    .Q(WX7787),
    .Q_t(WX7787_t)
  );


  xor2s3
  U821
  (
    .DIN1(n5283),
    .DIN1_t(n5283_t),
    .DIN2(n5463),
    .DIN2_t(n5463_t),
    .Q(n2781),
    .Q_t(n2781_t)
  );


  nor2s3
  U822
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n2782),
    .DIN2_t(n2782_t),
    .Q(WX7785),
    .Q_t(WX7785_t)
  );


  xor2s3
  U823
  (
    .DIN1(n5278),
    .DIN1_t(n5278_t),
    .DIN2(n5458),
    .DIN2_t(n5458_t),
    .Q(n2782),
    .Q_t(n2782_t)
  );


  nor2s3
  U824
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n2783),
    .DIN2_t(n2783_t),
    .Q(WX7783),
    .Q_t(WX7783_t)
  );


  xor2s3
  U825
  (
    .DIN1(n5273),
    .DIN1_t(n5273_t),
    .DIN2(n5453),
    .DIN2_t(n5453_t),
    .Q(n2783),
    .Q_t(n2783_t)
  );


  nor2s3
  U826
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n2784),
    .DIN2_t(n2784_t),
    .Q(WX7781),
    .Q_t(WX7781_t)
  );


  xor2s3
  U827
  (
    .DIN1(n5268),
    .DIN1_t(n5268_t),
    .DIN2(n5448),
    .DIN2_t(n5448_t),
    .Q(n2784),
    .Q_t(n2784_t)
  );


  nor2s3
  U828
  (
    .DIN1(n6485),
    .DIN1_t(n6485_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX778),
    .Q_t(WX778_t)
  );


  nor2s3
  U829
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n2785),
    .DIN2_t(n2785_t),
    .Q(WX7779),
    .Q_t(WX7779_t)
  );


  xor2s3
  U830
  (
    .DIN1(n5263),
    .DIN1_t(n5263_t),
    .DIN2(n5443),
    .DIN2_t(n5443_t),
    .Q(n2785),
    .Q_t(n2785_t)
  );


  nor2s3
  U831
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n2786),
    .DIN2_t(n2786_t),
    .Q(WX7777),
    .Q_t(WX7777_t)
  );


  xor2s3
  U832
  (
    .DIN1(n5258),
    .DIN1_t(n5258_t),
    .DIN2(n5438),
    .DIN2_t(n5438_t),
    .Q(n2786),
    .Q_t(n2786_t)
  );


  nor2s3
  U833
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2787),
    .DIN2_t(n2787_t),
    .Q(WX7775),
    .Q_t(WX7775_t)
  );


  xor2s3
  U834
  (
    .DIN1(n5253),
    .DIN1_t(n5253_t),
    .DIN2(n5433),
    .DIN2_t(n5433_t),
    .Q(n2787),
    .Q_t(n2787_t)
  );


  nor2s3
  U835
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2788),
    .DIN2_t(n2788_t),
    .Q(WX7773),
    .Q_t(WX7773_t)
  );


  xor2s3
  U836
  (
    .DIN1(n5248),
    .DIN1_t(n5248_t),
    .DIN2(n5428),
    .DIN2_t(n5428_t),
    .Q(n2788),
    .Q_t(n2788_t)
  );


  nor2s3
  U837
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2789),
    .DIN2_t(n2789_t),
    .Q(WX7771),
    .Q_t(WX7771_t)
  );


  xor2s3
  U838
  (
    .DIN1(n5243),
    .DIN1_t(n5243_t),
    .DIN2(n5423),
    .DIN2_t(n5423_t),
    .Q(n2789),
    .Q_t(n2789_t)
  );


  nor2s3
  U839
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2790),
    .DIN2_t(n2790_t),
    .Q(WX7769),
    .Q_t(WX7769_t)
  );


  xor2s3
  U840
  (
    .DIN1(n5238),
    .DIN1_t(n5238_t),
    .DIN2(n5418),
    .DIN2_t(n5418_t),
    .Q(n2790),
    .Q_t(n2790_t)
  );


  nor2s3
  U841
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2791),
    .DIN2_t(n2791_t),
    .Q(WX7767),
    .Q_t(WX7767_t)
  );


  xor2s3
  U842
  (
    .DIN1(n5233),
    .DIN1_t(n5233_t),
    .DIN2(n5413),
    .DIN2_t(n5413_t),
    .Q(n2791),
    .Q_t(n2791_t)
  );


  nor2s3
  U843
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2792),
    .DIN2_t(n2792_t),
    .Q(WX7765),
    .Q_t(WX7765_t)
  );


  xor2s3
  U844
  (
    .DIN1(n5228),
    .DIN1_t(n5228_t),
    .DIN2(n5408),
    .DIN2_t(n5408_t),
    .Q(n2792),
    .Q_t(n2792_t)
  );


  nor2s3
  U845
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2793),
    .DIN2_t(n2793_t),
    .Q(WX7763),
    .Q_t(WX7763_t)
  );


  xor2s3
  U846
  (
    .DIN1(n5223),
    .DIN1_t(n5223_t),
    .DIN2(n5403),
    .DIN2_t(n5403_t),
    .Q(n2793),
    .Q_t(n2793_t)
  );


  nor2s3
  U847
  (
    .DIN1(n2794),
    .DIN1_t(n2794_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX7761),
    .Q_t(WX7761_t)
  );


  xnr2s3
  U848
  (
    .DIN1(n5398),
    .DIN1_t(n5398_t),
    .DIN2(n2795),
    .DIN2_t(n2795_t),
    .Q(n2794),
    .Q_t(n2794_t)
  );


  xor2s3
  U849
  (
    .DIN1(n5218),
    .DIN1_t(n5218_t),
    .DIN2(n5298),
    .DIN2_t(n5298_t),
    .Q(n2795),
    .Q_t(n2795_t)
  );


  nor2s3
  U850
  (
    .DIN1(n6480),
    .DIN1_t(n6480_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX776),
    .Q_t(WX776_t)
  );


  nor2s3
  U851
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2796),
    .DIN2_t(n2796_t),
    .Q(WX7759),
    .Q_t(WX7759_t)
  );


  xor2s3
  U852
  (
    .DIN1(n5214),
    .DIN1_t(n5214_t),
    .DIN2(n3252),
    .DIN2_t(n3252_t),
    .Q(n2796),
    .Q_t(n2796_t)
  );


  nor2s3
  U853
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2797),
    .DIN2_t(n2797_t),
    .Q(WX7757),
    .Q_t(WX7757_t)
  );


  xor2s3
  U854
  (
    .DIN1(n5210),
    .DIN1_t(n5210_t),
    .DIN2(n3251),
    .DIN2_t(n3251_t),
    .Q(n2797),
    .Q_t(n2797_t)
  );


  nor2s3
  U855
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2798),
    .DIN2_t(n2798_t),
    .Q(WX7755),
    .Q_t(WX7755_t)
  );


  xor2s3
  U856
  (
    .DIN1(n5206),
    .DIN1_t(n5206_t),
    .DIN2(n3250),
    .DIN2_t(n3250_t),
    .Q(n2798),
    .Q_t(n2798_t)
  );


  nor2s3
  U857
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2799),
    .DIN2_t(n2799_t),
    .Q(WX7753),
    .Q_t(WX7753_t)
  );


  xor2s3
  U858
  (
    .DIN1(n5202),
    .DIN1_t(n5202_t),
    .DIN2(n3249),
    .DIN2_t(n3249_t),
    .Q(n2799),
    .Q_t(n2799_t)
  );


  nor2s3
  U859
  (
    .DIN1(n2800),
    .DIN1_t(n2800_t),
    .DIN2(n6746),
    .DIN2_t(n6746_t),
    .Q(WX7751),
    .Q_t(WX7751_t)
  );


  xnr2s3
  U860
  (
    .DIN1(n3248),
    .DIN1_t(n3248_t),
    .DIN2(n2801),
    .DIN2_t(n2801_t),
    .Q(n2800),
    .Q_t(n2800_t)
  );


  xor2s3
  U861
  (
    .DIN1(n5198),
    .DIN1_t(n5198_t),
    .DIN2(n5298),
    .DIN2_t(n5298_t),
    .Q(n2801),
    .Q_t(n2801_t)
  );


  nor2s3
  U862
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2802),
    .DIN2_t(n2802_t),
    .Q(WX7749),
    .Q_t(WX7749_t)
  );


  xor2s3
  U863
  (
    .DIN1(n5194),
    .DIN1_t(n5194_t),
    .DIN2(n3247),
    .DIN2_t(n3247_t),
    .Q(n2802),
    .Q_t(n2802_t)
  );


  nor2s3
  U864
  (
    .DIN1(n6801),
    .DIN1_t(n6801_t),
    .DIN2(n2803),
    .DIN2_t(n2803_t),
    .Q(WX7747),
    .Q_t(WX7747_t)
  );


  xor2s3
  U865
  (
    .DIN1(n5190),
    .DIN1_t(n5190_t),
    .DIN2(n3246),
    .DIN2_t(n3246_t),
    .Q(n2803),
    .Q_t(n2803_t)
  );


  nor2s3
  U866
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n2804),
    .DIN2_t(n2804_t),
    .Q(WX7745),
    .Q_t(WX7745_t)
  );


  xor2s3
  U867
  (
    .DIN1(n5186),
    .DIN1_t(n5186_t),
    .DIN2(n3245),
    .DIN2_t(n3245_t),
    .Q(n2804),
    .Q_t(n2804_t)
  );


  nor2s3
  U868
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n2805),
    .DIN2_t(n2805_t),
    .Q(WX7743),
    .Q_t(WX7743_t)
  );


  xor2s3
  U869
  (
    .DIN1(n5182),
    .DIN1_t(n5182_t),
    .DIN2(n3244),
    .DIN2_t(n3244_t),
    .Q(n2805),
    .Q_t(n2805_t)
  );


  nor2s3
  U870
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n2806),
    .DIN2_t(n2806_t),
    .Q(WX7741),
    .Q_t(WX7741_t)
  );


  xor2s3
  U871
  (
    .DIN1(n5178),
    .DIN1_t(n5178_t),
    .DIN2(n3243),
    .DIN2_t(n3243_t),
    .Q(n2806),
    .Q_t(n2806_t)
  );


  nor2s3
  U872
  (
    .DIN1(n6476),
    .DIN1_t(n6476_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX774),
    .Q_t(WX774_t)
  );


  nor2s3
  U873
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n2807),
    .DIN2_t(n2807_t),
    .Q(WX7739),
    .Q_t(WX7739_t)
  );


  xor2s3
  U874
  (
    .DIN1(n5174),
    .DIN1_t(n5174_t),
    .DIN2(n3242),
    .DIN2_t(n3242_t),
    .Q(n2807),
    .Q_t(n2807_t)
  );


  nor2s3
  U875
  (
    .DIN1(n2808),
    .DIN1_t(n2808_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX7737),
    .Q_t(WX7737_t)
  );


  xnr2s3
  U876
  (
    .DIN1(n3241),
    .DIN1_t(n3241_t),
    .DIN2(n2809),
    .DIN2_t(n2809_t),
    .Q(n2808),
    .Q_t(n2808_t)
  );


  xor2s3
  U877
  (
    .DIN1(n5170),
    .DIN1_t(n5170_t),
    .DIN2(n5298),
    .DIN2_t(n5298_t),
    .Q(n2809),
    .Q_t(n2809_t)
  );


  nor2s3
  U878
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n2810),
    .DIN2_t(n2810_t),
    .Q(WX7735),
    .Q_t(WX7735_t)
  );


  xor2s3
  U879
  (
    .DIN1(n5166),
    .DIN1_t(n5166_t),
    .DIN2(n3240),
    .DIN2_t(n3240_t),
    .Q(n2810),
    .Q_t(n2810_t)
  );


  nor2s3
  U880
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n2811),
    .DIN2_t(n2811_t),
    .Q(WX7733),
    .Q_t(WX7733_t)
  );


  xor2s3
  U881
  (
    .DIN1(n5162),
    .DIN1_t(n5162_t),
    .DIN2(n3239),
    .DIN2_t(n3239_t),
    .Q(n2811),
    .Q_t(n2811_t)
  );


  nor2s3
  U882
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n2812),
    .DIN2_t(n2812_t),
    .Q(WX7731),
    .Q_t(WX7731_t)
  );


  xor2s3
  U883
  (
    .DIN1(n5158),
    .DIN1_t(n5158_t),
    .DIN2(n3238),
    .DIN2_t(n3238_t),
    .Q(n2812),
    .Q_t(n2812_t)
  );


  nor2s3
  U884
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n2813),
    .DIN2_t(n2813_t),
    .Q(WX7729),
    .Q_t(WX7729_t)
  );


  xor2s3
  U885
  (
    .DIN1(n5298),
    .DIN1_t(n5298_t),
    .DIN2(n3237),
    .DIN2_t(n3237_t),
    .Q(n2813),
    .Q_t(n2813_t)
  );


  nor2s3
  U886
  (
    .DIN1(n6532),
    .DIN1_t(n6532_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX772),
    .Q_t(WX772_t)
  );


  nor2s3
  U887
  (
    .DIN1(n6553),
    .DIN1_t(n6553_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX770),
    .Q_t(WX770_t)
  );


  nor2s3
  U888
  (
    .DIN1(n6529),
    .DIN1_t(n6529_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX768),
    .Q_t(WX768_t)
  );


  nor2s3
  U889
  (
    .DIN1(n6435),
    .DIN1_t(n6435_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX766),
    .Q_t(WX766_t)
  );


  nor2s3
  U890
  (
    .DIN1(n6551),
    .DIN1_t(n6551_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX764),
    .Q_t(WX764_t)
  );


  nor2s3
  U891
  (
    .DIN1(n6550),
    .DIN1_t(n6550_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX762),
    .Q_t(WX762_t)
  );


  nor2s3
  U892
  (
    .DIN1(n6554),
    .DIN1_t(n6554_t),
    .DIN2(n6745),
    .DIN2_t(n6745_t),
    .Q(WX760),
    .Q_t(WX760_t)
  );


  nor2s3
  U893
  (
    .DIN1(n6560),
    .DIN1_t(n6560_t),
    .DIN2(n6750),
    .DIN2_t(n6750_t),
    .Q(WX758),
    .Q_t(WX758_t)
  );


  nor2s3
  U894
  (
    .DIN1(n6552),
    .DIN1_t(n6552_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX756),
    .Q_t(WX756_t)
  );


  nor2s3
  U895
  (
    .DIN1(n6556),
    .DIN1_t(n6556_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX754),
    .Q_t(WX754_t)
  );


  nor2s3
  U896
  (
    .DIN1(n6507),
    .DIN1_t(n6507_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX752),
    .Q_t(WX752_t)
  );


  nor2s3
  U897
  (
    .DIN1(n6557),
    .DIN1_t(n6557_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX750),
    .Q_t(WX750_t)
  );


  nor2s3
  U898
  (
    .DIN1(n6559),
    .DIN1_t(n6559_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX748),
    .Q_t(WX748_t)
  );


  nor2s3
  U899
  (
    .DIN1(n6555),
    .DIN1_t(n6555_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX746),
    .Q_t(WX746_t)
  );


  nor2s3
  U900
  (
    .DIN1(n6558),
    .DIN1_t(n6558_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX744),
    .Q_t(WX744_t)
  );


  nor2s3
  U901
  (
    .DIN1(n6526),
    .DIN1_t(n6526_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX742),
    .Q_t(WX742_t)
  );


  nor2s3
  U902
  (
    .DIN1(n6561),
    .DIN1_t(n6561_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX740),
    .Q_t(WX740_t)
  );


  nor2s3
  U903
  (
    .DIN1(n6509),
    .DIN1_t(n6509_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX738),
    .Q_t(WX738_t)
  );


  nor2s3
  U904
  (
    .DIN1(n5333),
    .DIN1_t(n5333_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX7363),
    .Q_t(WX7363_t)
  );


  nor2s3
  U905
  (
    .DIN1(n5337),
    .DIN1_t(n5337_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX7361),
    .Q_t(WX7361_t)
  );


  nor2s3
  U906
  (
    .DIN1(n6542),
    .DIN1_t(n6542_t),
    .DIN2(n6722),
    .DIN2_t(n6722_t),
    .Q(WX736),
    .Q_t(WX736_t)
  );


  nor2s3
  U907
  (
    .DIN1(n5341),
    .DIN1_t(n5341_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX7359),
    .Q_t(WX7359_t)
  );


  nor2s3
  U908
  (
    .DIN1(n5345),
    .DIN1_t(n5345_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX7357),
    .Q_t(WX7357_t)
  );


  nor2s3
  U909
  (
    .DIN1(n5349),
    .DIN1_t(n5349_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX7355),
    .Q_t(WX7355_t)
  );


  nor2s3
  U910
  (
    .DIN1(n5353),
    .DIN1_t(n5353_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX7353),
    .Q_t(WX7353_t)
  );


  nor2s3
  U911
  (
    .DIN1(n5357),
    .DIN1_t(n5357_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX7351),
    .Q_t(WX7351_t)
  );


  nor2s3
  U912
  (
    .DIN1(n5361),
    .DIN1_t(n5361_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX7349),
    .Q_t(WX7349_t)
  );


  nor2s3
  U913
  (
    .DIN1(n5365),
    .DIN1_t(n5365_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX7347),
    .Q_t(WX7347_t)
  );


  nor2s3
  U914
  (
    .DIN1(n5369),
    .DIN1_t(n5369_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX7345),
    .Q_t(WX7345_t)
  );


  nor2s3
  U915
  (
    .DIN1(n5373),
    .DIN1_t(n5373_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX7343),
    .Q_t(WX7343_t)
  );


  nor2s3
  U916
  (
    .DIN1(n5377),
    .DIN1_t(n5377_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX7341),
    .Q_t(WX7341_t)
  );


  nor2s3
  U917
  (
    .DIN1(n6490),
    .DIN1_t(n6490_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX734),
    .Q_t(WX734_t)
  );


  nor2s3
  U918
  (
    .DIN1(n5381),
    .DIN1_t(n5381_t),
    .DIN2(n6721),
    .DIN2_t(n6721_t),
    .Q(WX7339),
    .Q_t(WX7339_t)
  );


  nor2s3
  U919
  (
    .DIN1(n5385),
    .DIN1_t(n5385_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX7337),
    .Q_t(WX7337_t)
  );


  nor2s3
  U920
  (
    .DIN1(n5389),
    .DIN1_t(n5389_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX7335),
    .Q_t(WX7335_t)
  );


  nor2s3
  U921
  (
    .DIN1(n5393),
    .DIN1_t(n5393_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX7333),
    .Q_t(WX7333_t)
  );


  nor2s3
  U922
  (
    .DIN1(n5397),
    .DIN1_t(n5397_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX7331),
    .Q_t(WX7331_t)
  );


  nor2s3
  U923
  (
    .DIN1(n5402),
    .DIN1_t(n5402_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX7329),
    .Q_t(WX7329_t)
  );


  nor2s3
  U924
  (
    .DIN1(n5407),
    .DIN1_t(n5407_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX7327),
    .Q_t(WX7327_t)
  );


  nor2s3
  U925
  (
    .DIN1(n5412),
    .DIN1_t(n5412_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX7325),
    .Q_t(WX7325_t)
  );


  nor2s3
  U926
  (
    .DIN1(n5417),
    .DIN1_t(n5417_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX7323),
    .Q_t(WX7323_t)
  );


  nor2s3
  U927
  (
    .DIN1(n5422),
    .DIN1_t(n5422_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX7321),
    .Q_t(WX7321_t)
  );


  nor2s3
  U928
  (
    .DIN1(n6548),
    .DIN1_t(n6548_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX732),
    .Q_t(WX732_t)
  );


  nor2s3
  U929
  (
    .DIN1(n5427),
    .DIN1_t(n5427_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX7319),
    .Q_t(WX7319_t)
  );


  nor2s3
  U930
  (
    .DIN1(n5432),
    .DIN1_t(n5432_t),
    .DIN2(n6720),
    .DIN2_t(n6720_t),
    .Q(WX7317),
    .Q_t(WX7317_t)
  );


  nor2s3
  U931
  (
    .DIN1(n5437),
    .DIN1_t(n5437_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX7315),
    .Q_t(WX7315_t)
  );


  nor2s3
  U932
  (
    .DIN1(n5442),
    .DIN1_t(n5442_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX7313),
    .Q_t(WX7313_t)
  );


  nor2s3
  U933
  (
    .DIN1(n5447),
    .DIN1_t(n5447_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX7311),
    .Q_t(WX7311_t)
  );


  nor2s3
  U934
  (
    .DIN1(n5452),
    .DIN1_t(n5452_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX7309),
    .Q_t(WX7309_t)
  );


  nor2s3
  U935
  (
    .DIN1(n5457),
    .DIN1_t(n5457_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX7307),
    .Q_t(WX7307_t)
  );


  nor2s3
  U936
  (
    .DIN1(n5462),
    .DIN1_t(n5462_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX7305),
    .Q_t(WX7305_t)
  );


  nor2s3
  U937
  (
    .DIN1(n5467),
    .DIN1_t(n5467_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX7303),
    .Q_t(WX7303_t)
  );


  nor2s3
  U938
  (
    .DIN1(n5472),
    .DIN1_t(n5472_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX7301),
    .Q_t(WX7301_t)
  );


  nor2s3
  U939
  (
    .DIN1(n6521),
    .DIN1_t(n6521_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX730),
    .Q_t(WX730_t)
  );


  nor2s3
  U940
  (
    .DIN1(n5332),
    .DIN1_t(n5332_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX7299),
    .Q_t(WX7299_t)
  );


  nor2s3
  U941
  (
    .DIN1(n5336),
    .DIN1_t(n5336_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX7297),
    .Q_t(WX7297_t)
  );


  nor2s3
  U942
  (
    .DIN1(n5340),
    .DIN1_t(n5340_t),
    .DIN2(n6719),
    .DIN2_t(n6719_t),
    .Q(WX7295),
    .Q_t(WX7295_t)
  );


  nor2s3
  U943
  (
    .DIN1(n5344),
    .DIN1_t(n5344_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX7293),
    .Q_t(WX7293_t)
  );


  nor2s3
  U944
  (
    .DIN1(n5348),
    .DIN1_t(n5348_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX7291),
    .Q_t(WX7291_t)
  );


  nor2s3
  U945
  (
    .DIN1(n5352),
    .DIN1_t(n5352_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX7289),
    .Q_t(WX7289_t)
  );


  nor2s3
  U946
  (
    .DIN1(n5356),
    .DIN1_t(n5356_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX7287),
    .Q_t(WX7287_t)
  );


  nor2s3
  U947
  (
    .DIN1(n5360),
    .DIN1_t(n5360_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX7285),
    .Q_t(WX7285_t)
  );


  nor2s3
  U948
  (
    .DIN1(n5364),
    .DIN1_t(n5364_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX7283),
    .Q_t(WX7283_t)
  );


  nor2s3
  U949
  (
    .DIN1(n5368),
    .DIN1_t(n5368_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX7281),
    .Q_t(WX7281_t)
  );


  nor2s3
  U950
  (
    .DIN1(n6536),
    .DIN1_t(n6536_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX728),
    .Q_t(WX728_t)
  );


  nor2s3
  U951
  (
    .DIN1(n5372),
    .DIN1_t(n5372_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX7279),
    .Q_t(WX7279_t)
  );


  nor2s3
  U952
  (
    .DIN1(n5376),
    .DIN1_t(n5376_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX7277),
    .Q_t(WX7277_t)
  );


  nor2s3
  U953
  (
    .DIN1(n5380),
    .DIN1_t(n5380_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX7275),
    .Q_t(WX7275_t)
  );


  nor2s3
  U954
  (
    .DIN1(n5384),
    .DIN1_t(n5384_t),
    .DIN2(n6718),
    .DIN2_t(n6718_t),
    .Q(WX7273),
    .Q_t(WX7273_t)
  );


  nor2s3
  U955
  (
    .DIN1(n5388),
    .DIN1_t(n5388_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX7271),
    .Q_t(WX7271_t)
  );


  nor2s3
  U956
  (
    .DIN1(n5392),
    .DIN1_t(n5392_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX7269),
    .Q_t(WX7269_t)
  );


  and2s3
  U957
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5396),
    .DIN2_t(n5396_t),
    .Q(WX7267),
    .Q_t(WX7267_t)
  );


  and2s3
  U958
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5401),
    .DIN2_t(n5401_t),
    .Q(WX7265),
    .Q_t(WX7265_t)
  );


  and2s3
  U959
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5406),
    .DIN2_t(n5406_t),
    .Q(WX7263),
    .Q_t(WX7263_t)
  );


  and2s3
  U960
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5411),
    .DIN2_t(n5411_t),
    .Q(WX7261),
    .Q_t(WX7261_t)
  );


  nor2s3
  U961
  (
    .DIN1(n6515),
    .DIN1_t(n6515_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX726),
    .Q_t(WX726_t)
  );


  and2s3
  U962
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5416),
    .DIN2_t(n5416_t),
    .Q(WX7259),
    .Q_t(WX7259_t)
  );


  and2s3
  U963
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5421),
    .DIN2_t(n5421_t),
    .Q(WX7257),
    .Q_t(WX7257_t)
  );


  and2s3
  U964
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5426),
    .DIN2_t(n5426_t),
    .Q(WX7255),
    .Q_t(WX7255_t)
  );


  and2s3
  U965
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5431),
    .DIN2_t(n5431_t),
    .Q(WX7253),
    .Q_t(WX7253_t)
  );


  and2s3
  U966
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5436),
    .DIN2_t(n5436_t),
    .Q(WX7251),
    .Q_t(WX7251_t)
  );


  and2s3
  U967
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5441),
    .DIN2_t(n5441_t),
    .Q(WX7249),
    .Q_t(WX7249_t)
  );


  and2s3
  U968
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5446),
    .DIN2_t(n5446_t),
    .Q(WX7247),
    .Q_t(WX7247_t)
  );


  and2s3
  U969
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5451),
    .DIN2_t(n5451_t),
    .Q(WX7245),
    .Q_t(WX7245_t)
  );


  and2s3
  U970
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5456),
    .DIN2_t(n5456_t),
    .Q(WX7243),
    .Q_t(WX7243_t)
  );


  and2s3
  U971
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5461),
    .DIN2_t(n5461_t),
    .Q(WX7241),
    .Q_t(WX7241_t)
  );


  nor2s3
  U972
  (
    .DIN1(n6538),
    .DIN1_t(n6538_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX724),
    .Q_t(WX724_t)
  );


  and2s3
  U973
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5466),
    .DIN2_t(n5466_t),
    .Q(WX7239),
    .Q_t(WX7239_t)
  );


  and2s3
  U974
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5471),
    .DIN2_t(n5471_t),
    .Q(WX7237),
    .Q_t(WX7237_t)
  );


  and2s3
  U975
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5331),
    .DIN2_t(n5331_t),
    .Q(WX7235),
    .Q_t(WX7235_t)
  );


  and2s3
  U976
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5335),
    .DIN2_t(n5335_t),
    .Q(WX7233),
    .Q_t(WX7233_t)
  );


  and2s3
  U977
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5339),
    .DIN2_t(n5339_t),
    .Q(WX7231),
    .Q_t(WX7231_t)
  );


  and2s3
  U978
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5343),
    .DIN2_t(n5343_t),
    .Q(WX7229),
    .Q_t(WX7229_t)
  );


  and2s3
  U979
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5347),
    .DIN2_t(n5347_t),
    .Q(WX7227),
    .Q_t(WX7227_t)
  );


  and2s3
  U980
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5351),
    .DIN2_t(n5351_t),
    .Q(WX7225),
    .Q_t(WX7225_t)
  );


  and2s3
  U981
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5355),
    .DIN2_t(n5355_t),
    .Q(WX7223),
    .Q_t(WX7223_t)
  );


  and2s3
  U982
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5359),
    .DIN2_t(n5359_t),
    .Q(WX7221),
    .Q_t(WX7221_t)
  );


  nor2s3
  U983
  (
    .DIN1(n6540),
    .DIN1_t(n6540_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX722),
    .Q_t(WX722_t)
  );


  and2s3
  U984
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5363),
    .DIN2_t(n5363_t),
    .Q(WX7219),
    .Q_t(WX7219_t)
  );


  and2s3
  U985
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5367),
    .DIN2_t(n5367_t),
    .Q(WX7217),
    .Q_t(WX7217_t)
  );


  and2s3
  U986
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5371),
    .DIN2_t(n5371_t),
    .Q(WX7215),
    .Q_t(WX7215_t)
  );


  and2s3
  U987
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5375),
    .DIN2_t(n5375_t),
    .Q(WX7213),
    .Q_t(WX7213_t)
  );


  and2s3
  U988
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5379),
    .DIN2_t(n5379_t),
    .Q(WX7211),
    .Q_t(WX7211_t)
  );


  and2s3
  U989
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5383),
    .DIN2_t(n5383_t),
    .Q(WX7209),
    .Q_t(WX7209_t)
  );


  and2s3
  U990
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5387),
    .DIN2_t(n5387_t),
    .Q(WX7207),
    .Q_t(WX7207_t)
  );


  and2s3
  U991
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5391),
    .DIN2_t(n5391_t),
    .Q(WX7205),
    .Q_t(WX7205_t)
  );


  nor2s3
  U992
  (
    .DIN1(n5395),
    .DIN1_t(n5395_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX7203),
    .Q_t(WX7203_t)
  );


  nor2s3
  U993
  (
    .DIN1(n5400),
    .DIN1_t(n5400_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX7201),
    .Q_t(WX7201_t)
  );


  nor2s3
  U994
  (
    .DIN1(n6499),
    .DIN1_t(n6499_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX720),
    .Q_t(WX720_t)
  );


  nor2s3
  U995
  (
    .DIN1(n5405),
    .DIN1_t(n5405_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX7199),
    .Q_t(WX7199_t)
  );


  nor2s3
  U996
  (
    .DIN1(n5410),
    .DIN1_t(n5410_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX7197),
    .Q_t(WX7197_t)
  );


  nor2s3
  U997
  (
    .DIN1(n5415),
    .DIN1_t(n5415_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX7195),
    .Q_t(WX7195_t)
  );


  nor2s3
  U998
  (
    .DIN1(n5420),
    .DIN1_t(n5420_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX7193),
    .Q_t(WX7193_t)
  );


  nor2s3
  U999
  (
    .DIN1(n5425),
    .DIN1_t(n5425_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX7191),
    .Q_t(WX7191_t)
  );


  nor2s3
  U1000
  (
    .DIN1(n5430),
    .DIN1_t(n5430_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX7189),
    .Q_t(WX7189_t)
  );


  nor2s3
  U1001
  (
    .DIN1(n5435),
    .DIN1_t(n5435_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX7187),
    .Q_t(WX7187_t)
  );


  nor2s3
  U1002
  (
    .DIN1(n5440),
    .DIN1_t(n5440_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX7185),
    .Q_t(WX7185_t)
  );


  nor2s3
  U1003
  (
    .DIN1(n5445),
    .DIN1_t(n5445_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX7183),
    .Q_t(WX7183_t)
  );


  nor2s3
  U1004
  (
    .DIN1(n5450),
    .DIN1_t(n5450_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX7181),
    .Q_t(WX7181_t)
  );


  nor2s3
  U1005
  (
    .DIN1(n6543),
    .DIN1_t(n6543_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX718),
    .Q_t(WX718_t)
  );


  nor2s3
  U1006
  (
    .DIN1(n5455),
    .DIN1_t(n5455_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX7179),
    .Q_t(WX7179_t)
  );


  nor2s3
  U1007
  (
    .DIN1(n5460),
    .DIN1_t(n5460_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX7177),
    .Q_t(WX7177_t)
  );


  nor2s3
  U1008
  (
    .DIN1(n5465),
    .DIN1_t(n5465_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX7175),
    .Q_t(WX7175_t)
  );


  nor2s3
  U1009
  (
    .DIN1(n5470),
    .DIN1_t(n5470_t),
    .DIN2(n6716),
    .DIN2_t(n6716_t),
    .Q(WX7173),
    .Q_t(WX7173_t)
  );


  nnd4s2
  U1010
  (
    .DIN1(n2814),
    .DIN1_t(n2814_t),
    .DIN2(n2815),
    .DIN2_t(n2815_t),
    .DIN3(n2816),
    .DIN3_t(n2816_t),
    .DIN4(n2817),
    .DIN4_t(n2817_t),
    .Q(WX7171),
    .Q_t(WX7171_t)
  );


  nnd2s3
  U1011
  (
    .DIN1(n2545),
    .DIN1_t(n2545_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2817),
    .Q_t(n2817_t)
  );


  xor2s3
  U1012
  (
    .DIN1(n2818),
    .DIN1_t(n2818_t),
    .DIN2(n2819),
    .DIN2_t(n2819_t),
    .Q(n2545),
    .Q_t(n2545_t)
  );


  xor2s3
  U1013
  (
    .DIN1(n5155),
    .DIN1_t(n5155_t),
    .DIN2(n5156),
    .DIN2_t(n5156_t),
    .Q(n2819),
    .Q_t(n2819_t)
  );


  xnr2s3
  U1014
  (
    .DIN1(n3221),
    .DIN1_t(n3221_t),
    .DIN2(n5157),
    .DIN2_t(n5157_t),
    .Q(n2818),
    .Q_t(n2818_t)
  );


  nnd2s3
  U1015
  (
    .DIN1(n2820),
    .DIN1_t(n2820_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2816),
    .Q_t(n2816_t)
  );


  nnd2s3
  U1016
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1953),
    .DIN2_t(n1953_t),
    .Q(n2815),
    .Q_t(n2815_t)
  );


  nnd2s3
  U1017
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1952),
    .DIN2_t(n1952_t),
    .Q(n2814),
    .Q_t(n2814_t)
  );


  nnd4s2
  U1018
  (
    .DIN1(n2821),
    .DIN1_t(n2821_t),
    .DIN2(n2822),
    .DIN2_t(n2822_t),
    .DIN3(n2823),
    .DIN3_t(n2823_t),
    .DIN4(n2824),
    .DIN4_t(n2824_t),
    .Q(WX7169),
    .Q_t(WX7169_t)
  );


  nnd2s3
  U1019
  (
    .DIN1(n2552),
    .DIN1_t(n2552_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2824),
    .Q_t(n2824_t)
  );


  xor2s3
  U1020
  (
    .DIN1(n2825),
    .DIN1_t(n2825_t),
    .DIN2(n2826),
    .DIN2_t(n2826_t),
    .Q(n2552),
    .Q_t(n2552_t)
  );


  xor2s3
  U1021
  (
    .DIN1(n5159),
    .DIN1_t(n5159_t),
    .DIN2(n5160),
    .DIN2_t(n5160_t),
    .Q(n2826),
    .Q_t(n2826_t)
  );


  xnr2s3
  U1022
  (
    .DIN1(n3222),
    .DIN1_t(n3222_t),
    .DIN2(n5161),
    .DIN2_t(n5161_t),
    .Q(n2825),
    .Q_t(n2825_t)
  );


  nnd2s3
  U1023
  (
    .DIN1(n2827),
    .DIN1_t(n2827_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2823),
    .Q_t(n2823_t)
  );


  nnd2s3
  U1024
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1954),
    .DIN2_t(n1954_t),
    .Q(n2822),
    .Q_t(n2822_t)
  );


  nnd2s3
  U1025
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1951),
    .DIN2_t(n1951_t),
    .Q(n2821),
    .Q_t(n2821_t)
  );


  nnd4s2
  U1026
  (
    .DIN1(n2828),
    .DIN1_t(n2828_t),
    .DIN2(n2829),
    .DIN2_t(n2829_t),
    .DIN3(n2830),
    .DIN3_t(n2830_t),
    .DIN4(n2831),
    .DIN4_t(n2831_t),
    .Q(WX7167),
    .Q_t(WX7167_t)
  );


  nnd2s3
  U1027
  (
    .DIN1(n2559),
    .DIN1_t(n2559_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2831),
    .Q_t(n2831_t)
  );


  xor2s3
  U1028
  (
    .DIN1(n2832),
    .DIN1_t(n2832_t),
    .DIN2(n2833),
    .DIN2_t(n2833_t),
    .Q(n2559),
    .Q_t(n2559_t)
  );


  xor2s3
  U1029
  (
    .DIN1(n5163),
    .DIN1_t(n5163_t),
    .DIN2(n5164),
    .DIN2_t(n5164_t),
    .Q(n2833),
    .Q_t(n2833_t)
  );


  xnr2s3
  U1030
  (
    .DIN1(n3223),
    .DIN1_t(n3223_t),
    .DIN2(n5165),
    .DIN2_t(n5165_t),
    .Q(n2832),
    .Q_t(n2832_t)
  );


  nnd2s3
  U1031
  (
    .DIN1(n2834),
    .DIN1_t(n2834_t),
    .DIN2(n6662),
    .DIN2_t(n6662_t),
    .Q(n2830),
    .Q_t(n2830_t)
  );


  nnd2s3
  U1032
  (
    .DIN1(n6611),
    .DIN1_t(n6611_t),
    .DIN2(n1955),
    .DIN2_t(n1955_t),
    .Q(n2829),
    .Q_t(n2829_t)
  );


  nnd2s3
  U1033
  (
    .DIN1(n6580),
    .DIN1_t(n6580_t),
    .DIN2(n1950),
    .DIN2_t(n1950_t),
    .Q(n2828),
    .Q_t(n2828_t)
  );


  nnd4s2
  U1034
  (
    .DIN1(n2835),
    .DIN1_t(n2835_t),
    .DIN2(n2836),
    .DIN2_t(n2836_t),
    .DIN3(n2837),
    .DIN3_t(n2837_t),
    .DIN4(n2838),
    .DIN4_t(n2838_t),
    .Q(WX7165),
    .Q_t(WX7165_t)
  );


  nnd2s3
  U1035
  (
    .DIN1(n2566),
    .DIN1_t(n2566_t),
    .DIN2(n6631),
    .DIN2_t(n6631_t),
    .Q(n2838),
    .Q_t(n2838_t)
  );


  xor2s3
  U1036
  (
    .DIN1(n2839),
    .DIN1_t(n2839_t),
    .DIN2(n2840),
    .DIN2_t(n2840_t),
    .Q(n2566),
    .Q_t(n2566_t)
  );


  xor2s3
  U1037
  (
    .DIN1(n5167),
    .DIN1_t(n5167_t),
    .DIN2(n5168),
    .DIN2_t(n5168_t),
    .Q(n2840),
    .Q_t(n2840_t)
  );


  xnr2s3
  U1038
  (
    .DIN1(n3224),
    .DIN1_t(n3224_t),
    .DIN2(n5169),
    .DIN2_t(n5169_t),
    .Q(n2839),
    .Q_t(n2839_t)
  );


  nnd2s3
  U1039
  (
    .DIN1(n2841),
    .DIN1_t(n2841_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n2837),
    .Q_t(n2837_t)
  );


  nnd2s3
  U1040
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1956),
    .DIN2_t(n1956_t),
    .Q(n2836),
    .Q_t(n2836_t)
  );


  nnd2s3
  U1041
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1949),
    .DIN2_t(n1949_t),
    .Q(n2835),
    .Q_t(n2835_t)
  );


  nnd4s2
  U1042
  (
    .DIN1(n2842),
    .DIN1_t(n2842_t),
    .DIN2(n2843),
    .DIN2_t(n2843_t),
    .DIN3(n2844),
    .DIN3_t(n2844_t),
    .DIN4(n2845),
    .DIN4_t(n2845_t),
    .Q(WX7163),
    .Q_t(WX7163_t)
  );


  nnd2s3
  U1043
  (
    .DIN1(n2573),
    .DIN1_t(n2573_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n2845),
    .Q_t(n2845_t)
  );


  xor2s3
  U1044
  (
    .DIN1(n2846),
    .DIN1_t(n2846_t),
    .DIN2(n2847),
    .DIN2_t(n2847_t),
    .Q(n2573),
    .Q_t(n2573_t)
  );


  xor2s3
  U1045
  (
    .DIN1(n5171),
    .DIN1_t(n5171_t),
    .DIN2(n5172),
    .DIN2_t(n5172_t),
    .Q(n2847),
    .Q_t(n2847_t)
  );


  xnr2s3
  U1046
  (
    .DIN1(n3225),
    .DIN1_t(n3225_t),
    .DIN2(n5173),
    .DIN2_t(n5173_t),
    .Q(n2846),
    .Q_t(n2846_t)
  );


  nnd2s3
  U1047
  (
    .DIN1(n2848),
    .DIN1_t(n2848_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n2844),
    .Q_t(n2844_t)
  );


  nnd2s3
  U1048
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1957),
    .DIN2_t(n1957_t),
    .Q(n2843),
    .Q_t(n2843_t)
  );


  nnd2s3
  U1049
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1948),
    .DIN2_t(n1948_t),
    .Q(n2842),
    .Q_t(n2842_t)
  );


  nnd4s2
  U1050
  (
    .DIN1(n2849),
    .DIN1_t(n2849_t),
    .DIN2(n2850),
    .DIN2_t(n2850_t),
    .DIN3(n2851),
    .DIN3_t(n2851_t),
    .DIN4(n2852),
    .DIN4_t(n2852_t),
    .Q(WX7161),
    .Q_t(WX7161_t)
  );


  nnd2s3
  U1051
  (
    .DIN1(n2580),
    .DIN1_t(n2580_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n2852),
    .Q_t(n2852_t)
  );


  xor2s3
  U1052
  (
    .DIN1(n2853),
    .DIN1_t(n2853_t),
    .DIN2(n2854),
    .DIN2_t(n2854_t),
    .Q(n2580),
    .Q_t(n2580_t)
  );


  xor2s3
  U1053
  (
    .DIN1(n5175),
    .DIN1_t(n5175_t),
    .DIN2(n5176),
    .DIN2_t(n5176_t),
    .Q(n2854),
    .Q_t(n2854_t)
  );


  xnr2s3
  U1054
  (
    .DIN1(n3226),
    .DIN1_t(n3226_t),
    .DIN2(n5177),
    .DIN2_t(n5177_t),
    .Q(n2853),
    .Q_t(n2853_t)
  );


  nnd2s3
  U1055
  (
    .DIN1(n2855),
    .DIN1_t(n2855_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n2851),
    .Q_t(n2851_t)
  );


  nnd2s3
  U1056
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1958),
    .DIN2_t(n1958_t),
    .Q(n2850),
    .Q_t(n2850_t)
  );


  nnd2s3
  U1057
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1947),
    .DIN2_t(n1947_t),
    .Q(n2849),
    .Q_t(n2849_t)
  );


  nor2s3
  U1058
  (
    .DIN1(n6545),
    .DIN1_t(n6545_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX716),
    .Q_t(WX716_t)
  );


  nnd4s2
  U1059
  (
    .DIN1(n2856),
    .DIN1_t(n2856_t),
    .DIN2(n2857),
    .DIN2_t(n2857_t),
    .DIN3(n2858),
    .DIN3_t(n2858_t),
    .DIN4(n2859),
    .DIN4_t(n2859_t),
    .Q(WX7159),
    .Q_t(WX7159_t)
  );


  nnd2s3
  U1060
  (
    .DIN1(n2587),
    .DIN1_t(n2587_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n2859),
    .Q_t(n2859_t)
  );


  xor2s3
  U1061
  (
    .DIN1(n2860),
    .DIN1_t(n2860_t),
    .DIN2(n2861),
    .DIN2_t(n2861_t),
    .Q(n2587),
    .Q_t(n2587_t)
  );


  xor2s3
  U1062
  (
    .DIN1(n5179),
    .DIN1_t(n5179_t),
    .DIN2(n5180),
    .DIN2_t(n5180_t),
    .Q(n2861),
    .Q_t(n2861_t)
  );


  xnr2s3
  U1063
  (
    .DIN1(n3227),
    .DIN1_t(n3227_t),
    .DIN2(n5181),
    .DIN2_t(n5181_t),
    .Q(n2860),
    .Q_t(n2860_t)
  );


  nnd2s3
  U1064
  (
    .DIN1(n2862),
    .DIN1_t(n2862_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n2858),
    .Q_t(n2858_t)
  );


  nnd2s3
  U1065
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1959),
    .DIN2_t(n1959_t),
    .Q(n2857),
    .Q_t(n2857_t)
  );


  nnd2s3
  U1066
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1946),
    .DIN2_t(n1946_t),
    .Q(n2856),
    .Q_t(n2856_t)
  );


  nnd4s2
  U1067
  (
    .DIN1(n2863),
    .DIN1_t(n2863_t),
    .DIN2(n2864),
    .DIN2_t(n2864_t),
    .DIN3(n2865),
    .DIN3_t(n2865_t),
    .DIN4(n2866),
    .DIN4_t(n2866_t),
    .Q(WX7157),
    .Q_t(WX7157_t)
  );


  nnd2s3
  U1068
  (
    .DIN1(n2594),
    .DIN1_t(n2594_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n2866),
    .Q_t(n2866_t)
  );


  xor2s3
  U1069
  (
    .DIN1(n2867),
    .DIN1_t(n2867_t),
    .DIN2(n2868),
    .DIN2_t(n2868_t),
    .Q(n2594),
    .Q_t(n2594_t)
  );


  xor2s3
  U1070
  (
    .DIN1(n5183),
    .DIN1_t(n5183_t),
    .DIN2(n5184),
    .DIN2_t(n5184_t),
    .Q(n2868),
    .Q_t(n2868_t)
  );


  xnr2s3
  U1071
  (
    .DIN1(n3228),
    .DIN1_t(n3228_t),
    .DIN2(n5185),
    .DIN2_t(n5185_t),
    .Q(n2867),
    .Q_t(n2867_t)
  );


  nnd2s3
  U1072
  (
    .DIN1(n2869),
    .DIN1_t(n2869_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n2865),
    .Q_t(n2865_t)
  );


  nnd2s3
  U1073
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1960),
    .DIN2_t(n1960_t),
    .Q(n2864),
    .Q_t(n2864_t)
  );


  nnd2s3
  U1074
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1945),
    .DIN2_t(n1945_t),
    .Q(n2863),
    .Q_t(n2863_t)
  );


  nnd4s2
  U1075
  (
    .DIN1(n2870),
    .DIN1_t(n2870_t),
    .DIN2(n2871),
    .DIN2_t(n2871_t),
    .DIN3(n2872),
    .DIN3_t(n2872_t),
    .DIN4(n2873),
    .DIN4_t(n2873_t),
    .Q(WX7155),
    .Q_t(WX7155_t)
  );


  nnd2s3
  U1076
  (
    .DIN1(n2601),
    .DIN1_t(n2601_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n2873),
    .Q_t(n2873_t)
  );


  xor2s3
  U1077
  (
    .DIN1(n2874),
    .DIN1_t(n2874_t),
    .DIN2(n2875),
    .DIN2_t(n2875_t),
    .Q(n2601),
    .Q_t(n2601_t)
  );


  xor2s3
  U1078
  (
    .DIN1(n5187),
    .DIN1_t(n5187_t),
    .DIN2(n5188),
    .DIN2_t(n5188_t),
    .Q(n2875),
    .Q_t(n2875_t)
  );


  xnr2s3
  U1079
  (
    .DIN1(n3229),
    .DIN1_t(n3229_t),
    .DIN2(n5189),
    .DIN2_t(n5189_t),
    .Q(n2874),
    .Q_t(n2874_t)
  );


  nnd2s3
  U1080
  (
    .DIN1(n2876),
    .DIN1_t(n2876_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n2872),
    .Q_t(n2872_t)
  );


  nnd2s3
  U1081
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1961),
    .DIN2_t(n1961_t),
    .Q(n2871),
    .Q_t(n2871_t)
  );


  nnd2s3
  U1082
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1944),
    .DIN2_t(n1944_t),
    .Q(n2870),
    .Q_t(n2870_t)
  );


  nnd4s2
  U1083
  (
    .DIN1(n2877),
    .DIN1_t(n2877_t),
    .DIN2(n2878),
    .DIN2_t(n2878_t),
    .DIN3(n2879),
    .DIN3_t(n2879_t),
    .DIN4(n2880),
    .DIN4_t(n2880_t),
    .Q(WX7153),
    .Q_t(WX7153_t)
  );


  nnd2s3
  U1084
  (
    .DIN1(n2608),
    .DIN1_t(n2608_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n2880),
    .Q_t(n2880_t)
  );


  xor2s3
  U1085
  (
    .DIN1(n2881),
    .DIN1_t(n2881_t),
    .DIN2(n2882),
    .DIN2_t(n2882_t),
    .Q(n2608),
    .Q_t(n2608_t)
  );


  xor2s3
  U1086
  (
    .DIN1(n5191),
    .DIN1_t(n5191_t),
    .DIN2(n5192),
    .DIN2_t(n5192_t),
    .Q(n2882),
    .Q_t(n2882_t)
  );


  xnr2s3
  U1087
  (
    .DIN1(n3230),
    .DIN1_t(n3230_t),
    .DIN2(n5193),
    .DIN2_t(n5193_t),
    .Q(n2881),
    .Q_t(n2881_t)
  );


  nnd2s3
  U1088
  (
    .DIN1(n2883),
    .DIN1_t(n2883_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n2879),
    .Q_t(n2879_t)
  );


  nnd2s3
  U1089
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1962),
    .DIN2_t(n1962_t),
    .Q(n2878),
    .Q_t(n2878_t)
  );


  nnd2s3
  U1090
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1943),
    .DIN2_t(n1943_t),
    .Q(n2877),
    .Q_t(n2877_t)
  );


  nnd4s2
  U1091
  (
    .DIN1(n2884),
    .DIN1_t(n2884_t),
    .DIN2(n2885),
    .DIN2_t(n2885_t),
    .DIN3(n2886),
    .DIN3_t(n2886_t),
    .DIN4(n2887),
    .DIN4_t(n2887_t),
    .Q(WX7151),
    .Q_t(WX7151_t)
  );


  nnd2s3
  U1092
  (
    .DIN1(n2615),
    .DIN1_t(n2615_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n2887),
    .Q_t(n2887_t)
  );


  xor2s3
  U1093
  (
    .DIN1(n2888),
    .DIN1_t(n2888_t),
    .DIN2(n2889),
    .DIN2_t(n2889_t),
    .Q(n2615),
    .Q_t(n2615_t)
  );


  xor2s3
  U1094
  (
    .DIN1(n5195),
    .DIN1_t(n5195_t),
    .DIN2(n5196),
    .DIN2_t(n5196_t),
    .Q(n2889),
    .Q_t(n2889_t)
  );


  xnr2s3
  U1095
  (
    .DIN1(n3231),
    .DIN1_t(n3231_t),
    .DIN2(n5197),
    .DIN2_t(n5197_t),
    .Q(n2888),
    .Q_t(n2888_t)
  );


  nnd2s3
  U1096
  (
    .DIN1(n2890),
    .DIN1_t(n2890_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n2886),
    .Q_t(n2886_t)
  );


  nnd2s3
  U1097
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1963),
    .DIN2_t(n1963_t),
    .Q(n2885),
    .Q_t(n2885_t)
  );


  nnd2s3
  U1098
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1942),
    .DIN2_t(n1942_t),
    .Q(n2884),
    .Q_t(n2884_t)
  );


  nnd4s2
  U1099
  (
    .DIN1(n2891),
    .DIN1_t(n2891_t),
    .DIN2(n2892),
    .DIN2_t(n2892_t),
    .DIN3(n2893),
    .DIN3_t(n2893_t),
    .DIN4(n2894),
    .DIN4_t(n2894_t),
    .Q(WX7149),
    .Q_t(WX7149_t)
  );


  nnd2s3
  U1100
  (
    .DIN1(n2622),
    .DIN1_t(n2622_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n2894),
    .Q_t(n2894_t)
  );


  xor2s3
  U1101
  (
    .DIN1(n2895),
    .DIN1_t(n2895_t),
    .DIN2(n2896),
    .DIN2_t(n2896_t),
    .Q(n2622),
    .Q_t(n2622_t)
  );


  xor2s3
  U1102
  (
    .DIN1(n5199),
    .DIN1_t(n5199_t),
    .DIN2(n5200),
    .DIN2_t(n5200_t),
    .Q(n2896),
    .Q_t(n2896_t)
  );


  xnr2s3
  U1103
  (
    .DIN1(n3232),
    .DIN1_t(n3232_t),
    .DIN2(n5201),
    .DIN2_t(n5201_t),
    .Q(n2895),
    .Q_t(n2895_t)
  );


  nnd2s3
  U1104
  (
    .DIN1(n2897),
    .DIN1_t(n2897_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n2893),
    .Q_t(n2893_t)
  );


  nnd2s3
  U1105
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1964),
    .DIN2_t(n1964_t),
    .Q(n2892),
    .Q_t(n2892_t)
  );


  nnd2s3
  U1106
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1941),
    .DIN2_t(n1941_t),
    .Q(n2891),
    .Q_t(n2891_t)
  );


  nnd4s2
  U1107
  (
    .DIN1(n2898),
    .DIN1_t(n2898_t),
    .DIN2(n2899),
    .DIN2_t(n2899_t),
    .DIN3(n2900),
    .DIN3_t(n2900_t),
    .DIN4(n2901),
    .DIN4_t(n2901_t),
    .Q(WX7147),
    .Q_t(WX7147_t)
  );


  nnd2s3
  U1108
  (
    .DIN1(n2629),
    .DIN1_t(n2629_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n2901),
    .Q_t(n2901_t)
  );


  xor2s3
  U1109
  (
    .DIN1(n2902),
    .DIN1_t(n2902_t),
    .DIN2(n2903),
    .DIN2_t(n2903_t),
    .Q(n2629),
    .Q_t(n2629_t)
  );


  xor2s3
  U1110
  (
    .DIN1(n5203),
    .DIN1_t(n5203_t),
    .DIN2(n5204),
    .DIN2_t(n5204_t),
    .Q(n2903),
    .Q_t(n2903_t)
  );


  xnr2s3
  U1111
  (
    .DIN1(n3233),
    .DIN1_t(n3233_t),
    .DIN2(n5205),
    .DIN2_t(n5205_t),
    .Q(n2902),
    .Q_t(n2902_t)
  );


  nnd2s3
  U1112
  (
    .DIN1(n2904),
    .DIN1_t(n2904_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n2900),
    .Q_t(n2900_t)
  );


  nnd2s3
  U1113
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1965),
    .DIN2_t(n1965_t),
    .Q(n2899),
    .Q_t(n2899_t)
  );


  nnd2s3
  U1114
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1940),
    .DIN2_t(n1940_t),
    .Q(n2898),
    .Q_t(n2898_t)
  );


  nnd4s2
  U1115
  (
    .DIN1(n2905),
    .DIN1_t(n2905_t),
    .DIN2(n2906),
    .DIN2_t(n2906_t),
    .DIN3(n2907),
    .DIN3_t(n2907_t),
    .DIN4(n2908),
    .DIN4_t(n2908_t),
    .Q(WX7145),
    .Q_t(WX7145_t)
  );


  nnd2s3
  U1116
  (
    .DIN1(n2636),
    .DIN1_t(n2636_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n2908),
    .Q_t(n2908_t)
  );


  xor2s3
  U1117
  (
    .DIN1(n2909),
    .DIN1_t(n2909_t),
    .DIN2(n2910),
    .DIN2_t(n2910_t),
    .Q(n2636),
    .Q_t(n2636_t)
  );


  xor2s3
  U1118
  (
    .DIN1(n5207),
    .DIN1_t(n5207_t),
    .DIN2(n5208),
    .DIN2_t(n5208_t),
    .Q(n2910),
    .Q_t(n2910_t)
  );


  xnr2s3
  U1119
  (
    .DIN1(n3234),
    .DIN1_t(n3234_t),
    .DIN2(n5209),
    .DIN2_t(n5209_t),
    .Q(n2909),
    .Q_t(n2909_t)
  );


  nnd2s3
  U1120
  (
    .DIN1(n2911),
    .DIN1_t(n2911_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n2907),
    .Q_t(n2907_t)
  );


  nnd2s3
  U1121
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1966),
    .DIN2_t(n1966_t),
    .Q(n2906),
    .Q_t(n2906_t)
  );


  nnd2s3
  U1122
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1939),
    .DIN2_t(n1939_t),
    .Q(n2905),
    .Q_t(n2905_t)
  );


  nnd4s2
  U1123
  (
    .DIN1(n2912),
    .DIN1_t(n2912_t),
    .DIN2(n2913),
    .DIN2_t(n2913_t),
    .DIN3(n2914),
    .DIN3_t(n2914_t),
    .DIN4(n2915),
    .DIN4_t(n2915_t),
    .Q(WX7143),
    .Q_t(WX7143_t)
  );


  nnd2s3
  U1124
  (
    .DIN1(n2643),
    .DIN1_t(n2643_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n2915),
    .Q_t(n2915_t)
  );


  xor2s3
  U1125
  (
    .DIN1(n2916),
    .DIN1_t(n2916_t),
    .DIN2(n2917),
    .DIN2_t(n2917_t),
    .Q(n2643),
    .Q_t(n2643_t)
  );


  xor2s3
  U1126
  (
    .DIN1(n5211),
    .DIN1_t(n5211_t),
    .DIN2(n5212),
    .DIN2_t(n5212_t),
    .Q(n2917),
    .Q_t(n2917_t)
  );


  xnr2s3
  U1127
  (
    .DIN1(n3235),
    .DIN1_t(n3235_t),
    .DIN2(n5213),
    .DIN2_t(n5213_t),
    .Q(n2916),
    .Q_t(n2916_t)
  );


  nnd2s3
  U1128
  (
    .DIN1(n2918),
    .DIN1_t(n2918_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n2914),
    .Q_t(n2914_t)
  );


  nnd2s3
  U1129
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1967),
    .DIN2_t(n1967_t),
    .Q(n2913),
    .Q_t(n2913_t)
  );


  nnd2s3
  U1130
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1938),
    .DIN2_t(n1938_t),
    .Q(n2912),
    .Q_t(n2912_t)
  );


  nnd4s2
  U1131
  (
    .DIN1(n2919),
    .DIN1_t(n2919_t),
    .DIN2(n2920),
    .DIN2_t(n2920_t),
    .DIN3(n2921),
    .DIN3_t(n2921_t),
    .DIN4(n2922),
    .DIN4_t(n2922_t),
    .Q(WX7141),
    .Q_t(WX7141_t)
  );


  nnd2s3
  U1132
  (
    .DIN1(n2650),
    .DIN1_t(n2650_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n2922),
    .Q_t(n2922_t)
  );


  xor2s3
  U1133
  (
    .DIN1(n2923),
    .DIN1_t(n2923_t),
    .DIN2(n2924),
    .DIN2_t(n2924_t),
    .Q(n2650),
    .Q_t(n2650_t)
  );


  xor2s3
  U1134
  (
    .DIN1(n5215),
    .DIN1_t(n5215_t),
    .DIN2(n5216),
    .DIN2_t(n5216_t),
    .Q(n2924),
    .Q_t(n2924_t)
  );


  xnr2s3
  U1135
  (
    .DIN1(n3236),
    .DIN1_t(n3236_t),
    .DIN2(n5217),
    .DIN2_t(n5217_t),
    .Q(n2923),
    .Q_t(n2923_t)
  );


  nnd2s3
  U1136
  (
    .DIN1(n2925),
    .DIN1_t(n2925_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n2921),
    .Q_t(n2921_t)
  );


  nnd2s3
  U1137
  (
    .DIN1(n6610),
    .DIN1_t(n6610_t),
    .DIN2(n1968),
    .DIN2_t(n1968_t),
    .Q(n2920),
    .Q_t(n2920_t)
  );


  nnd2s3
  U1138
  (
    .DIN1(n6579),
    .DIN1_t(n6579_t),
    .DIN2(n1937),
    .DIN2_t(n1937_t),
    .Q(n2919),
    .Q_t(n2919_t)
  );


  nor2s3
  U1139
  (
    .DIN1(n6546),
    .DIN1_t(n6546_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX714),
    .Q_t(WX714_t)
  );


  nnd4s2
  U1140
  (
    .DIN1(n2926),
    .DIN1_t(n2926_t),
    .DIN2(n2927),
    .DIN2_t(n2927_t),
    .DIN3(n2928),
    .DIN3_t(n2928_t),
    .DIN4(n2929),
    .DIN4_t(n2929_t),
    .Q(WX7139),
    .Q_t(WX7139_t)
  );


  nnd2s3
  U1141
  (
    .DIN1(n2658),
    .DIN1_t(n2658_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n2929),
    .Q_t(n2929_t)
  );


  xor2s3
  U1142
  (
    .DIN1(n2930),
    .DIN1_t(n2930_t),
    .DIN2(n2931),
    .DIN2_t(n2931_t),
    .Q(n2658),
    .Q_t(n2658_t)
  );


  xor2s3
  U1143
  (
    .DIN1(n5221),
    .DIN1_t(n5221_t),
    .DIN2(n2932),
    .DIN2_t(n2932_t),
    .Q(n2931),
    .Q_t(n2931_t)
  );


  xor2s3
  U1144
  (
    .DIN1(n5219),
    .DIN1_t(n5219_t),
    .DIN2(n5220),
    .DIN2_t(n5220_t),
    .Q(n2932),
    .Q_t(n2932_t)
  );


  xor2s3
  U1145
  (
    .DIN1(n5222),
    .DIN1_t(n5222_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2930),
    .Q_t(n2930_t)
  );


  nnd2s3
  U1146
  (
    .DIN1(n2933),
    .DIN1_t(n2933_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n2928),
    .Q_t(n2928_t)
  );


  nnd2s3
  U1147
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1969),
    .DIN2_t(n1969_t),
    .Q(n2927),
    .Q_t(n2927_t)
  );


  nnd2s3
  U1148
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1936),
    .DIN2_t(n1936_t),
    .Q(n2926),
    .Q_t(n2926_t)
  );


  nnd4s2
  U1149
  (
    .DIN1(n2934),
    .DIN1_t(n2934_t),
    .DIN2(n2935),
    .DIN2_t(n2935_t),
    .DIN3(n2936),
    .DIN3_t(n2936_t),
    .DIN4(n2937),
    .DIN4_t(n2937_t),
    .Q(WX7137),
    .Q_t(WX7137_t)
  );


  nnd2s3
  U1150
  (
    .DIN1(n2666),
    .DIN1_t(n2666_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n2937),
    .Q_t(n2937_t)
  );


  xor2s3
  U1151
  (
    .DIN1(n2938),
    .DIN1_t(n2938_t),
    .DIN2(n2939),
    .DIN2_t(n2939_t),
    .Q(n2666),
    .Q_t(n2666_t)
  );


  xor2s3
  U1152
  (
    .DIN1(n5226),
    .DIN1_t(n5226_t),
    .DIN2(n2940),
    .DIN2_t(n2940_t),
    .Q(n2939),
    .Q_t(n2939_t)
  );


  xor2s3
  U1153
  (
    .DIN1(n5224),
    .DIN1_t(n5224_t),
    .DIN2(n5225),
    .DIN2_t(n5225_t),
    .Q(n2940),
    .Q_t(n2940_t)
  );


  xor2s3
  U1154
  (
    .DIN1(n5227),
    .DIN1_t(n5227_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2938),
    .Q_t(n2938_t)
  );


  nnd2s3
  U1155
  (
    .DIN1(n2941),
    .DIN1_t(n2941_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n2936),
    .Q_t(n2936_t)
  );


  nnd2s3
  U1156
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1970),
    .DIN2_t(n1970_t),
    .Q(n2935),
    .Q_t(n2935_t)
  );


  nnd2s3
  U1157
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1935),
    .DIN2_t(n1935_t),
    .Q(n2934),
    .Q_t(n2934_t)
  );


  nnd4s2
  U1158
  (
    .DIN1(n2942),
    .DIN1_t(n2942_t),
    .DIN2(n2943),
    .DIN2_t(n2943_t),
    .DIN3(n2944),
    .DIN3_t(n2944_t),
    .DIN4(n2945),
    .DIN4_t(n2945_t),
    .Q(WX7135),
    .Q_t(WX7135_t)
  );


  nnd2s3
  U1159
  (
    .DIN1(n2674),
    .DIN1_t(n2674_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n2945),
    .Q_t(n2945_t)
  );


  xor2s3
  U1160
  (
    .DIN1(n2946),
    .DIN1_t(n2946_t),
    .DIN2(n2947),
    .DIN2_t(n2947_t),
    .Q(n2674),
    .Q_t(n2674_t)
  );


  xor2s3
  U1161
  (
    .DIN1(n5231),
    .DIN1_t(n5231_t),
    .DIN2(n2948),
    .DIN2_t(n2948_t),
    .Q(n2947),
    .Q_t(n2947_t)
  );


  xor2s3
  U1162
  (
    .DIN1(n5229),
    .DIN1_t(n5229_t),
    .DIN2(n5230),
    .DIN2_t(n5230_t),
    .Q(n2948),
    .Q_t(n2948_t)
  );


  xor2s3
  U1163
  (
    .DIN1(n5232),
    .DIN1_t(n5232_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2946),
    .Q_t(n2946_t)
  );


  nnd2s3
  U1164
  (
    .DIN1(n2949),
    .DIN1_t(n2949_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n2944),
    .Q_t(n2944_t)
  );


  nnd2s3
  U1165
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1971),
    .DIN2_t(n1971_t),
    .Q(n2943),
    .Q_t(n2943_t)
  );


  nnd2s3
  U1166
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1934),
    .DIN2_t(n1934_t),
    .Q(n2942),
    .Q_t(n2942_t)
  );


  nnd4s2
  U1167
  (
    .DIN1(n2950),
    .DIN1_t(n2950_t),
    .DIN2(n2951),
    .DIN2_t(n2951_t),
    .DIN3(n2952),
    .DIN3_t(n2952_t),
    .DIN4(n2953),
    .DIN4_t(n2953_t),
    .Q(WX7133),
    .Q_t(WX7133_t)
  );


  nnd2s3
  U1168
  (
    .DIN1(n2682),
    .DIN1_t(n2682_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n2953),
    .Q_t(n2953_t)
  );


  xor2s3
  U1169
  (
    .DIN1(n2954),
    .DIN1_t(n2954_t),
    .DIN2(n2955),
    .DIN2_t(n2955_t),
    .Q(n2682),
    .Q_t(n2682_t)
  );


  xor2s3
  U1170
  (
    .DIN1(n5236),
    .DIN1_t(n5236_t),
    .DIN2(n2956),
    .DIN2_t(n2956_t),
    .Q(n2955),
    .Q_t(n2955_t)
  );


  xor2s3
  U1171
  (
    .DIN1(n5234),
    .DIN1_t(n5234_t),
    .DIN2(n5235),
    .DIN2_t(n5235_t),
    .Q(n2956),
    .Q_t(n2956_t)
  );


  xor2s3
  U1172
  (
    .DIN1(n5237),
    .DIN1_t(n5237_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2954),
    .Q_t(n2954_t)
  );


  nnd2s3
  U1173
  (
    .DIN1(n2957),
    .DIN1_t(n2957_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n2952),
    .Q_t(n2952_t)
  );


  nnd2s3
  U1174
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1972),
    .DIN2_t(n1972_t),
    .Q(n2951),
    .Q_t(n2951_t)
  );


  nnd2s3
  U1175
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1933),
    .DIN2_t(n1933_t),
    .Q(n2950),
    .Q_t(n2950_t)
  );


  nnd4s2
  U1176
  (
    .DIN1(n2958),
    .DIN1_t(n2958_t),
    .DIN2(n2959),
    .DIN2_t(n2959_t),
    .DIN3(n2960),
    .DIN3_t(n2960_t),
    .DIN4(n2961),
    .DIN4_t(n2961_t),
    .Q(WX7131),
    .Q_t(WX7131_t)
  );


  nnd2s3
  U1177
  (
    .DIN1(n2690),
    .DIN1_t(n2690_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n2961),
    .Q_t(n2961_t)
  );


  xor2s3
  U1178
  (
    .DIN1(n2962),
    .DIN1_t(n2962_t),
    .DIN2(n2963),
    .DIN2_t(n2963_t),
    .Q(n2690),
    .Q_t(n2690_t)
  );


  xor2s3
  U1179
  (
    .DIN1(n5241),
    .DIN1_t(n5241_t),
    .DIN2(n2964),
    .DIN2_t(n2964_t),
    .Q(n2963),
    .Q_t(n2963_t)
  );


  xor2s3
  U1180
  (
    .DIN1(n5239),
    .DIN1_t(n5239_t),
    .DIN2(n5240),
    .DIN2_t(n5240_t),
    .Q(n2964),
    .Q_t(n2964_t)
  );


  xor2s3
  U1181
  (
    .DIN1(n5242),
    .DIN1_t(n5242_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2962),
    .Q_t(n2962_t)
  );


  nnd2s3
  U1182
  (
    .DIN1(n2965),
    .DIN1_t(n2965_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n2960),
    .Q_t(n2960_t)
  );


  nnd2s3
  U1183
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1973),
    .DIN2_t(n1973_t),
    .Q(n2959),
    .Q_t(n2959_t)
  );


  nnd2s3
  U1184
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1932),
    .DIN2_t(n1932_t),
    .Q(n2958),
    .Q_t(n2958_t)
  );


  nnd4s2
  U1185
  (
    .DIN1(n2966),
    .DIN1_t(n2966_t),
    .DIN2(n2967),
    .DIN2_t(n2967_t),
    .DIN3(n2968),
    .DIN3_t(n2968_t),
    .DIN4(n2969),
    .DIN4_t(n2969_t),
    .Q(WX7129),
    .Q_t(WX7129_t)
  );


  nnd2s3
  U1186
  (
    .DIN1(n2698),
    .DIN1_t(n2698_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n2969),
    .Q_t(n2969_t)
  );


  xor2s3
  U1187
  (
    .DIN1(n2970),
    .DIN1_t(n2970_t),
    .DIN2(n2971),
    .DIN2_t(n2971_t),
    .Q(n2698),
    .Q_t(n2698_t)
  );


  xor2s3
  U1188
  (
    .DIN1(n5246),
    .DIN1_t(n5246_t),
    .DIN2(n2972),
    .DIN2_t(n2972_t),
    .Q(n2971),
    .Q_t(n2971_t)
  );


  xor2s3
  U1189
  (
    .DIN1(n5244),
    .DIN1_t(n5244_t),
    .DIN2(n5245),
    .DIN2_t(n5245_t),
    .Q(n2972),
    .Q_t(n2972_t)
  );


  xor2s3
  U1190
  (
    .DIN1(n5247),
    .DIN1_t(n5247_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2970),
    .Q_t(n2970_t)
  );


  nnd2s3
  U1191
  (
    .DIN1(n2973),
    .DIN1_t(n2973_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n2968),
    .Q_t(n2968_t)
  );


  nnd2s3
  U1192
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1974),
    .DIN2_t(n1974_t),
    .Q(n2967),
    .Q_t(n2967_t)
  );


  nnd2s3
  U1193
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1931),
    .DIN2_t(n1931_t),
    .Q(n2966),
    .Q_t(n2966_t)
  );


  nnd4s2
  U1194
  (
    .DIN1(n2974),
    .DIN1_t(n2974_t),
    .DIN2(n2975),
    .DIN2_t(n2975_t),
    .DIN3(n2976),
    .DIN3_t(n2976_t),
    .DIN4(n2977),
    .DIN4_t(n2977_t),
    .Q(WX7127),
    .Q_t(WX7127_t)
  );


  nnd2s3
  U1195
  (
    .DIN1(n2706),
    .DIN1_t(n2706_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n2977),
    .Q_t(n2977_t)
  );


  xor2s3
  U1196
  (
    .DIN1(n2978),
    .DIN1_t(n2978_t),
    .DIN2(n2979),
    .DIN2_t(n2979_t),
    .Q(n2706),
    .Q_t(n2706_t)
  );


  xor2s3
  U1197
  (
    .DIN1(n5251),
    .DIN1_t(n5251_t),
    .DIN2(n2980),
    .DIN2_t(n2980_t),
    .Q(n2979),
    .Q_t(n2979_t)
  );


  xor2s3
  U1198
  (
    .DIN1(n5249),
    .DIN1_t(n5249_t),
    .DIN2(n5250),
    .DIN2_t(n5250_t),
    .Q(n2980),
    .Q_t(n2980_t)
  );


  xor2s3
  U1199
  (
    .DIN1(n5252),
    .DIN1_t(n5252_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2978),
    .Q_t(n2978_t)
  );


  nnd2s3
  U1200
  (
    .DIN1(n2981),
    .DIN1_t(n2981_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n2976),
    .Q_t(n2976_t)
  );


  nnd2s3
  U1201
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1975),
    .DIN2_t(n1975_t),
    .Q(n2975),
    .Q_t(n2975_t)
  );


  nnd2s3
  U1202
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1930),
    .DIN2_t(n1930_t),
    .Q(n2974),
    .Q_t(n2974_t)
  );


  nnd4s2
  U1203
  (
    .DIN1(n2982),
    .DIN1_t(n2982_t),
    .DIN2(n2983),
    .DIN2_t(n2983_t),
    .DIN3(n2984),
    .DIN3_t(n2984_t),
    .DIN4(n2985),
    .DIN4_t(n2985_t),
    .Q(WX7125),
    .Q_t(WX7125_t)
  );


  nnd2s3
  U1204
  (
    .DIN1(n2714),
    .DIN1_t(n2714_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n2985),
    .Q_t(n2985_t)
  );


  xor2s3
  U1205
  (
    .DIN1(n2986),
    .DIN1_t(n2986_t),
    .DIN2(n2987),
    .DIN2_t(n2987_t),
    .Q(n2714),
    .Q_t(n2714_t)
  );


  xor2s3
  U1206
  (
    .DIN1(n5256),
    .DIN1_t(n5256_t),
    .DIN2(n2988),
    .DIN2_t(n2988_t),
    .Q(n2987),
    .Q_t(n2987_t)
  );


  xor2s3
  U1207
  (
    .DIN1(n5254),
    .DIN1_t(n5254_t),
    .DIN2(n5255),
    .DIN2_t(n5255_t),
    .Q(n2988),
    .Q_t(n2988_t)
  );


  xor2s3
  U1208
  (
    .DIN1(n5257),
    .DIN1_t(n5257_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2986),
    .Q_t(n2986_t)
  );


  nnd2s3
  U1209
  (
    .DIN1(n2989),
    .DIN1_t(n2989_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n2984),
    .Q_t(n2984_t)
  );


  nnd2s3
  U1210
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1976),
    .DIN2_t(n1976_t),
    .Q(n2983),
    .Q_t(n2983_t)
  );


  nnd2s3
  U1211
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1929),
    .DIN2_t(n1929_t),
    .Q(n2982),
    .Q_t(n2982_t)
  );


  nnd4s2
  U1212
  (
    .DIN1(n2990),
    .DIN1_t(n2990_t),
    .DIN2(n2991),
    .DIN2_t(n2991_t),
    .DIN3(n2992),
    .DIN3_t(n2992_t),
    .DIN4(n2993),
    .DIN4_t(n2993_t),
    .Q(WX7123),
    .Q_t(WX7123_t)
  );


  nnd2s3
  U1213
  (
    .DIN1(n2722),
    .DIN1_t(n2722_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n2993),
    .Q_t(n2993_t)
  );


  xor2s3
  U1214
  (
    .DIN1(n2994),
    .DIN1_t(n2994_t),
    .DIN2(n2995),
    .DIN2_t(n2995_t),
    .Q(n2722),
    .Q_t(n2722_t)
  );


  xor2s3
  U1215
  (
    .DIN1(n5261),
    .DIN1_t(n5261_t),
    .DIN2(n2996),
    .DIN2_t(n2996_t),
    .Q(n2995),
    .Q_t(n2995_t)
  );


  xor2s3
  U1216
  (
    .DIN1(n5259),
    .DIN1_t(n5259_t),
    .DIN2(n5260),
    .DIN2_t(n5260_t),
    .Q(n2996),
    .Q_t(n2996_t)
  );


  xor2s3
  U1217
  (
    .DIN1(n5262),
    .DIN1_t(n5262_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n2994),
    .Q_t(n2994_t)
  );


  nnd2s3
  U1218
  (
    .DIN1(n2997),
    .DIN1_t(n2997_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n2992),
    .Q_t(n2992_t)
  );


  nnd2s3
  U1219
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1977),
    .DIN2_t(n1977_t),
    .Q(n2991),
    .Q_t(n2991_t)
  );


  nnd2s3
  U1220
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1928),
    .DIN2_t(n1928_t),
    .Q(n2990),
    .Q_t(n2990_t)
  );


  nnd4s2
  U1221
  (
    .DIN1(n2998),
    .DIN1_t(n2998_t),
    .DIN2(n2999),
    .DIN2_t(n2999_t),
    .DIN3(n3000),
    .DIN3_t(n3000_t),
    .DIN4(n3001),
    .DIN4_t(n3001_t),
    .Q(WX7121),
    .Q_t(WX7121_t)
  );


  nnd2s3
  U1222
  (
    .DIN1(n2730),
    .DIN1_t(n2730_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n3001),
    .Q_t(n3001_t)
  );


  xor2s3
  U1223
  (
    .DIN1(n3002),
    .DIN1_t(n3002_t),
    .DIN2(n3003),
    .DIN2_t(n3003_t),
    .Q(n2730),
    .Q_t(n2730_t)
  );


  xor2s3
  U1224
  (
    .DIN1(n5266),
    .DIN1_t(n5266_t),
    .DIN2(n3004),
    .DIN2_t(n3004_t),
    .Q(n3003),
    .Q_t(n3003_t)
  );


  xor2s3
  U1225
  (
    .DIN1(n5264),
    .DIN1_t(n5264_t),
    .DIN2(n5265),
    .DIN2_t(n5265_t),
    .Q(n3004),
    .Q_t(n3004_t)
  );


  xor2s3
  U1226
  (
    .DIN1(n5267),
    .DIN1_t(n5267_t),
    .DIN2(n6688),
    .DIN2_t(n6688_t),
    .Q(n3002),
    .Q_t(n3002_t)
  );


  nnd2s3
  U1227
  (
    .DIN1(n3005),
    .DIN1_t(n3005_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n3000),
    .Q_t(n3000_t)
  );


  nnd2s3
  U1228
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1978),
    .DIN2_t(n1978_t),
    .Q(n2999),
    .Q_t(n2999_t)
  );


  nnd2s3
  U1229
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1927),
    .DIN2_t(n1927_t),
    .Q(n2998),
    .Q_t(n2998_t)
  );


  nor2s3
  U1230
  (
    .DIN1(n6481),
    .DIN1_t(n6481_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX712),
    .Q_t(WX712_t)
  );


  nnd4s2
  U1231
  (
    .DIN1(n3006),
    .DIN1_t(n3006_t),
    .DIN2(n3007),
    .DIN2_t(n3007_t),
    .DIN3(n3008),
    .DIN3_t(n3008_t),
    .DIN4(n3009),
    .DIN4_t(n3009_t),
    .Q(WX7119),
    .Q_t(WX7119_t)
  );


  nnd2s3
  U1232
  (
    .DIN1(n2738),
    .DIN1_t(n2738_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n3009),
    .Q_t(n3009_t)
  );


  xor2s3
  U1233
  (
    .DIN1(n3010),
    .DIN1_t(n3010_t),
    .DIN2(n3011),
    .DIN2_t(n3011_t),
    .Q(n2738),
    .Q_t(n2738_t)
  );


  xor2s3
  U1234
  (
    .DIN1(n5271),
    .DIN1_t(n5271_t),
    .DIN2(n3012),
    .DIN2_t(n3012_t),
    .Q(n3011),
    .Q_t(n3011_t)
  );


  xor2s3
  U1235
  (
    .DIN1(n5269),
    .DIN1_t(n5269_t),
    .DIN2(n5270),
    .DIN2_t(n5270_t),
    .Q(n3012),
    .Q_t(n3012_t)
  );


  xor2s3
  U1236
  (
    .DIN1(n5272),
    .DIN1_t(n5272_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3010),
    .Q_t(n3010_t)
  );


  nnd2s3
  U1237
  (
    .DIN1(n3013),
    .DIN1_t(n3013_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n3008),
    .Q_t(n3008_t)
  );


  nnd2s3
  U1238
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1979),
    .DIN2_t(n1979_t),
    .Q(n3007),
    .Q_t(n3007_t)
  );


  nnd2s3
  U1239
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1926),
    .DIN2_t(n1926_t),
    .Q(n3006),
    .Q_t(n3006_t)
  );


  nnd4s2
  U1240
  (
    .DIN1(n3014),
    .DIN1_t(n3014_t),
    .DIN2(n3015),
    .DIN2_t(n3015_t),
    .DIN3(n3016),
    .DIN3_t(n3016_t),
    .DIN4(n3017),
    .DIN4_t(n3017_t),
    .Q(WX7117),
    .Q_t(WX7117_t)
  );


  nnd2s3
  U1241
  (
    .DIN1(n2746),
    .DIN1_t(n2746_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n3017),
    .Q_t(n3017_t)
  );


  xor2s3
  U1242
  (
    .DIN1(n3018),
    .DIN1_t(n3018_t),
    .DIN2(n3019),
    .DIN2_t(n3019_t),
    .Q(n2746),
    .Q_t(n2746_t)
  );


  xor2s3
  U1243
  (
    .DIN1(n5276),
    .DIN1_t(n5276_t),
    .DIN2(n3020),
    .DIN2_t(n3020_t),
    .Q(n3019),
    .Q_t(n3019_t)
  );


  xor2s3
  U1244
  (
    .DIN1(n5274),
    .DIN1_t(n5274_t),
    .DIN2(n5275),
    .DIN2_t(n5275_t),
    .Q(n3020),
    .Q_t(n3020_t)
  );


  xor2s3
  U1245
  (
    .DIN1(n5277),
    .DIN1_t(n5277_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3018),
    .Q_t(n3018_t)
  );


  nnd2s3
  U1246
  (
    .DIN1(n3021),
    .DIN1_t(n3021_t),
    .DIN2(n6660),
    .DIN2_t(n6660_t),
    .Q(n3016),
    .Q_t(n3016_t)
  );


  nnd2s3
  U1247
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1980),
    .DIN2_t(n1980_t),
    .Q(n3015),
    .Q_t(n3015_t)
  );


  nnd2s3
  U1248
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1925),
    .DIN2_t(n1925_t),
    .Q(n3014),
    .Q_t(n3014_t)
  );


  nnd4s2
  U1249
  (
    .DIN1(n3022),
    .DIN1_t(n3022_t),
    .DIN2(n3023),
    .DIN2_t(n3023_t),
    .DIN3(n3024),
    .DIN3_t(n3024_t),
    .DIN4(n3025),
    .DIN4_t(n3025_t),
    .Q(WX7115),
    .Q_t(WX7115_t)
  );


  nnd2s3
  U1250
  (
    .DIN1(n2754),
    .DIN1_t(n2754_t),
    .DIN2(n6629),
    .DIN2_t(n6629_t),
    .Q(n3025),
    .Q_t(n3025_t)
  );


  xor2s3
  U1251
  (
    .DIN1(n3026),
    .DIN1_t(n3026_t),
    .DIN2(n3027),
    .DIN2_t(n3027_t),
    .Q(n2754),
    .Q_t(n2754_t)
  );


  xor2s3
  U1252
  (
    .DIN1(n5281),
    .DIN1_t(n5281_t),
    .DIN2(n3028),
    .DIN2_t(n3028_t),
    .Q(n3027),
    .Q_t(n3027_t)
  );


  xor2s3
  U1253
  (
    .DIN1(n5279),
    .DIN1_t(n5279_t),
    .DIN2(n5280),
    .DIN2_t(n5280_t),
    .Q(n3028),
    .Q_t(n3028_t)
  );


  xor2s3
  U1254
  (
    .DIN1(n5282),
    .DIN1_t(n5282_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3026),
    .Q_t(n3026_t)
  );


  nnd2s3
  U1255
  (
    .DIN1(n3029),
    .DIN1_t(n3029_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3024),
    .Q_t(n3024_t)
  );


  nnd2s3
  U1256
  (
    .DIN1(n6609),
    .DIN1_t(n6609_t),
    .DIN2(n1981),
    .DIN2_t(n1981_t),
    .Q(n3023),
    .Q_t(n3023_t)
  );


  nnd2s3
  U1257
  (
    .DIN1(n6578),
    .DIN1_t(n6578_t),
    .DIN2(n1924),
    .DIN2_t(n1924_t),
    .Q(n3022),
    .Q_t(n3022_t)
  );


  nnd4s2
  U1258
  (
    .DIN1(n3030),
    .DIN1_t(n3030_t),
    .DIN2(n3031),
    .DIN2_t(n3031_t),
    .DIN3(n3032),
    .DIN3_t(n3032_t),
    .DIN4(n3033),
    .DIN4_t(n3033_t),
    .Q(WX7113),
    .Q_t(WX7113_t)
  );


  nnd2s3
  U1259
  (
    .DIN1(n2762),
    .DIN1_t(n2762_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3033),
    .Q_t(n3033_t)
  );


  xor2s3
  U1260
  (
    .DIN1(n3034),
    .DIN1_t(n3034_t),
    .DIN2(n3035),
    .DIN2_t(n3035_t),
    .Q(n2762),
    .Q_t(n2762_t)
  );


  xor2s3
  U1261
  (
    .DIN1(n5286),
    .DIN1_t(n5286_t),
    .DIN2(n3036),
    .DIN2_t(n3036_t),
    .Q(n3035),
    .Q_t(n3035_t)
  );


  xor2s3
  U1262
  (
    .DIN1(n5284),
    .DIN1_t(n5284_t),
    .DIN2(n5285),
    .DIN2_t(n5285_t),
    .Q(n3036),
    .Q_t(n3036_t)
  );


  xor2s3
  U1263
  (
    .DIN1(n5287),
    .DIN1_t(n5287_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3034),
    .Q_t(n3034_t)
  );


  nnd2s3
  U1264
  (
    .DIN1(n3037),
    .DIN1_t(n3037_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3032),
    .Q_t(n3032_t)
  );


  nnd2s3
  U1265
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n1982),
    .DIN2_t(n1982_t),
    .Q(n3031),
    .Q_t(n3031_t)
  );


  nnd2s3
  U1266
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n1923),
    .DIN2_t(n1923_t),
    .Q(n3030),
    .Q_t(n3030_t)
  );


  nnd4s2
  U1267
  (
    .DIN1(n3038),
    .DIN1_t(n3038_t),
    .DIN2(n3039),
    .DIN2_t(n3039_t),
    .DIN3(n3040),
    .DIN3_t(n3040_t),
    .DIN4(n3041),
    .DIN4_t(n3041_t),
    .Q(WX7111),
    .Q_t(WX7111_t)
  );


  nnd2s3
  U1268
  (
    .DIN1(n2770),
    .DIN1_t(n2770_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3041),
    .Q_t(n3041_t)
  );


  xor2s3
  U1269
  (
    .DIN1(n3042),
    .DIN1_t(n3042_t),
    .DIN2(n3043),
    .DIN2_t(n3043_t),
    .Q(n2770),
    .Q_t(n2770_t)
  );


  xor2s3
  U1270
  (
    .DIN1(n5291),
    .DIN1_t(n5291_t),
    .DIN2(n3044),
    .DIN2_t(n3044_t),
    .Q(n3043),
    .Q_t(n3043_t)
  );


  xor2s3
  U1271
  (
    .DIN1(n5289),
    .DIN1_t(n5289_t),
    .DIN2(n5290),
    .DIN2_t(n5290_t),
    .Q(n3044),
    .Q_t(n3044_t)
  );


  xor2s3
  U1272
  (
    .DIN1(n5292),
    .DIN1_t(n5292_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3042),
    .Q_t(n3042_t)
  );


  nnd2s3
  U1273
  (
    .DIN1(n3045),
    .DIN1_t(n3045_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3040),
    .Q_t(n3040_t)
  );


  nnd2s3
  U1274
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n1983),
    .DIN2_t(n1983_t),
    .Q(n3039),
    .Q_t(n3039_t)
  );


  nnd2s3
  U1275
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n1922),
    .DIN2_t(n1922_t),
    .Q(n3038),
    .Q_t(n3038_t)
  );


  nnd4s2
  U1276
  (
    .DIN1(n3046),
    .DIN1_t(n3046_t),
    .DIN2(n3047),
    .DIN2_t(n3047_t),
    .DIN3(n3048),
    .DIN3_t(n3048_t),
    .DIN4(n3049),
    .DIN4_t(n3049_t),
    .Q(WX7109),
    .Q_t(WX7109_t)
  );


  nnd2s3
  U1277
  (
    .DIN1(n2778),
    .DIN1_t(n2778_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3049),
    .Q_t(n3049_t)
  );


  xor2s3
  U1278
  (
    .DIN1(n3050),
    .DIN1_t(n3050_t),
    .DIN2(n3051),
    .DIN2_t(n3051_t),
    .Q(n2778),
    .Q_t(n2778_t)
  );


  xor2s3
  U1279
  (
    .DIN1(n5296),
    .DIN1_t(n5296_t),
    .DIN2(n3052),
    .DIN2_t(n3052_t),
    .Q(n3051),
    .Q_t(n3051_t)
  );


  xor2s3
  U1280
  (
    .DIN1(n5294),
    .DIN1_t(n5294_t),
    .DIN2(n5295),
    .DIN2_t(n5295_t),
    .Q(n3052),
    .Q_t(n3052_t)
  );


  xor2s3
  U1281
  (
    .DIN1(n5297),
    .DIN1_t(n5297_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3050),
    .Q_t(n3050_t)
  );


  nnd2s3
  U1282
  (
    .DIN1(n3053),
    .DIN1_t(n3053_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3048),
    .Q_t(n3048_t)
  );


  nnd2s3
  U1283
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n1984),
    .DIN2_t(n1984_t),
    .Q(n3047),
    .Q_t(n3047_t)
  );


  nnd2s3
  U1284
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n1921),
    .DIN2_t(n1921_t),
    .Q(n3046),
    .Q_t(n3046_t)
  );


  nor2s3
  U1285
  (
    .DIN1(n6549),
    .DIN1_t(n6549_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX710),
    .Q_t(WX710_t)
  );


  nor2s3
  U1286
  (
    .DIN1(n6533),
    .DIN1_t(n6533_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX708),
    .Q_t(WX708_t)
  );


  nnd4s2
  U1287
  (
    .DIN1(n3054),
    .DIN1_t(n3054_t),
    .DIN2(n3055),
    .DIN2_t(n3055_t),
    .DIN3(n3056),
    .DIN3_t(n3056_t),
    .DIN4(n3057),
    .DIN4_t(n3057_t),
    .Q(WX706),
    .Q_t(WX706_t)
  );


  nnd2s3
  U1288
  (
    .DIN1(n3058),
    .DIN1_t(n3058_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3057),
    .Q_t(n3057_t)
  );


  nnd2s3
  U1289
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n2273),
    .DIN2_t(n2273_t),
    .Q(n3056),
    .Q_t(n3056_t)
  );


  nnd2s3
  U1290
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n2272),
    .DIN2_t(n2272_t),
    .Q(n3055),
    .Q_t(n3055_t)
  );


  nnd2s3
  U1291
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3059),
    .DIN2_t(n3059_t),
    .Q(n3054),
    .Q_t(n3054_t)
  );


  nnd4s2
  U1292
  (
    .DIN1(n3060),
    .DIN1_t(n3060_t),
    .DIN2(n3061),
    .DIN2_t(n3061_t),
    .DIN3(n3062),
    .DIN3_t(n3062_t),
    .DIN4(n3063),
    .DIN4_t(n3063_t),
    .Q(WX704),
    .Q_t(WX704_t)
  );


  nnd2s3
  U1293
  (
    .DIN1(n3064),
    .DIN1_t(n3064_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3063),
    .Q_t(n3063_t)
  );


  nnd2s3
  U1294
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n2274),
    .DIN2_t(n2274_t),
    .Q(n3062),
    .Q_t(n3062_t)
  );


  nnd2s3
  U1295
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n2271),
    .DIN2_t(n2271_t),
    .Q(n3061),
    .Q_t(n3061_t)
  );


  nnd2s3
  U1296
  (
    .DIN1(n6658),
    .DIN1_t(n6658_t),
    .DIN2(n3065),
    .DIN2_t(n3065_t),
    .Q(n3060),
    .Q_t(n3060_t)
  );


  nnd4s2
  U1297
  (
    .DIN1(n3066),
    .DIN1_t(n3066_t),
    .DIN2(n3067),
    .DIN2_t(n3067_t),
    .DIN3(n3068),
    .DIN3_t(n3068_t),
    .DIN4(n3069),
    .DIN4_t(n3069_t),
    .Q(WX702),
    .Q_t(WX702_t)
  );


  nnd2s3
  U1298
  (
    .DIN1(n3070),
    .DIN1_t(n3070_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3069),
    .Q_t(n3069_t)
  );


  nnd2s3
  U1299
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n2275),
    .DIN2_t(n2275_t),
    .Q(n3068),
    .Q_t(n3068_t)
  );


  nnd2s3
  U1300
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n2270),
    .DIN2_t(n2270_t),
    .Q(n3067),
    .Q_t(n3067_t)
  );


  nnd2s3
  U1301
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3071),
    .DIN2_t(n3071_t),
    .Q(n3066),
    .Q_t(n3066_t)
  );


  nor2s3
  U1302
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n1984),
    .DIN2_t(n1984_t),
    .Q(WX7011),
    .Q_t(WX7011_t)
  );


  nor2s3
  U1303
  (
    .DIN1(n5300),
    .DIN1_t(n5300_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX7009),
    .Q_t(WX7009_t)
  );


  nor2s3
  U1304
  (
    .DIN1(n5301),
    .DIN1_t(n5301_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX7007),
    .Q_t(WX7007_t)
  );


  nor2s3
  U1305
  (
    .DIN1(n5302),
    .DIN1_t(n5302_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX7005),
    .Q_t(WX7005_t)
  );


  nor2s3
  U1306
  (
    .DIN1(n5303),
    .DIN1_t(n5303_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX7003),
    .Q_t(WX7003_t)
  );


  nor2s3
  U1307
  (
    .DIN1(n5304),
    .DIN1_t(n5304_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX7001),
    .Q_t(WX7001_t)
  );


  nnd4s2
  U1308
  (
    .DIN1(n3072),
    .DIN1_t(n3072_t),
    .DIN2(n3073),
    .DIN2_t(n3073_t),
    .DIN3(n3074),
    .DIN3_t(n3074_t),
    .DIN4(n3075),
    .DIN4_t(n3075_t),
    .Q(WX700),
    .Q_t(WX700_t)
  );


  nnd2s3
  U1309
  (
    .DIN1(n3076),
    .DIN1_t(n3076_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3075),
    .Q_t(n3075_t)
  );


  nnd2s3
  U1310
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n2276),
    .DIN2_t(n2276_t),
    .Q(n3074),
    .Q_t(n3074_t)
  );


  nnd2s3
  U1311
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n2269),
    .DIN2_t(n2269_t),
    .Q(n3073),
    .Q_t(n3073_t)
  );


  nnd2s3
  U1312
  (
    .DIN1(n6658),
    .DIN1_t(n6658_t),
    .DIN2(n3077),
    .DIN2_t(n3077_t),
    .Q(n3072),
    .Q_t(n3072_t)
  );


  nor2s3
  U1313
  (
    .DIN1(n5305),
    .DIN1_t(n5305_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX6999),
    .Q_t(WX6999_t)
  );


  nor2s3
  U1314
  (
    .DIN1(n5306),
    .DIN1_t(n5306_t),
    .DIN2(n6715),
    .DIN2_t(n6715_t),
    .Q(WX6997),
    .Q_t(WX6997_t)
  );


  nor2s3
  U1315
  (
    .DIN1(n5307),
    .DIN1_t(n5307_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6995),
    .Q_t(WX6995_t)
  );


  nor2s3
  U1316
  (
    .DIN1(n5308),
    .DIN1_t(n5308_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6993),
    .Q_t(WX6993_t)
  );


  nor2s3
  U1317
  (
    .DIN1(n5309),
    .DIN1_t(n5309_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6991),
    .Q_t(WX6991_t)
  );


  nor2s3
  U1318
  (
    .DIN1(n5310),
    .DIN1_t(n5310_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6989),
    .Q_t(WX6989_t)
  );


  nor2s3
  U1319
  (
    .DIN1(n5311),
    .DIN1_t(n5311_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6987),
    .Q_t(WX6987_t)
  );


  nor2s3
  U1320
  (
    .DIN1(n5312),
    .DIN1_t(n5312_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6985),
    .Q_t(WX6985_t)
  );


  nor2s3
  U1321
  (
    .DIN1(n5313),
    .DIN1_t(n5313_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6983),
    .Q_t(WX6983_t)
  );


  nor2s3
  U1322
  (
    .DIN1(n5314),
    .DIN1_t(n5314_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6981),
    .Q_t(WX6981_t)
  );


  nnd4s2
  U1323
  (
    .DIN1(n3078),
    .DIN1_t(n3078_t),
    .DIN2(n3079),
    .DIN2_t(n3079_t),
    .DIN3(n3080),
    .DIN3_t(n3080_t),
    .DIN4(n3081),
    .DIN4_t(n3081_t),
    .Q(WX698),
    .Q_t(WX698_t)
  );


  nnd2s3
  U1324
  (
    .DIN1(n3082),
    .DIN1_t(n3082_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3081),
    .Q_t(n3081_t)
  );


  nnd2s3
  U1325
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n2277),
    .DIN2_t(n2277_t),
    .Q(n3080),
    .Q_t(n3080_t)
  );


  nnd2s3
  U1326
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n2268),
    .DIN2_t(n2268_t),
    .Q(n3079),
    .Q_t(n3079_t)
  );


  nnd2s3
  U1327
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3083),
    .DIN2_t(n3083_t),
    .Q(n3078),
    .Q_t(n3078_t)
  );


  nor2s3
  U1328
  (
    .DIN1(n5315),
    .DIN1_t(n5315_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6979),
    .Q_t(WX6979_t)
  );


  nor2s3
  U1329
  (
    .DIN1(n5316),
    .DIN1_t(n5316_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6977),
    .Q_t(WX6977_t)
  );


  nor2s3
  U1330
  (
    .DIN1(n5317),
    .DIN1_t(n5317_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6975),
    .Q_t(WX6975_t)
  );


  nor2s3
  U1331
  (
    .DIN1(n5318),
    .DIN1_t(n5318_t),
    .DIN2(n6714),
    .DIN2_t(n6714_t),
    .Q(WX6973),
    .Q_t(WX6973_t)
  );


  nor2s3
  U1332
  (
    .DIN1(n5319),
    .DIN1_t(n5319_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6971),
    .Q_t(WX6971_t)
  );


  nor2s3
  U1333
  (
    .DIN1(n5320),
    .DIN1_t(n5320_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6969),
    .Q_t(WX6969_t)
  );


  nor2s3
  U1334
  (
    .DIN1(n5321),
    .DIN1_t(n5321_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6967),
    .Q_t(WX6967_t)
  );


  nor2s3
  U1335
  (
    .DIN1(n5322),
    .DIN1_t(n5322_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6965),
    .Q_t(WX6965_t)
  );


  nor2s3
  U1336
  (
    .DIN1(n5323),
    .DIN1_t(n5323_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6963),
    .Q_t(WX6963_t)
  );


  nor2s3
  U1337
  (
    .DIN1(n5324),
    .DIN1_t(n5324_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6961),
    .Q_t(WX6961_t)
  );


  nnd4s2
  U1338
  (
    .DIN1(n3084),
    .DIN1_t(n3084_t),
    .DIN2(n3085),
    .DIN2_t(n3085_t),
    .DIN3(n3086),
    .DIN3_t(n3086_t),
    .DIN4(n3087),
    .DIN4_t(n3087_t),
    .Q(WX696),
    .Q_t(WX696_t)
  );


  nnd2s3
  U1339
  (
    .DIN1(n3088),
    .DIN1_t(n3088_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3087),
    .Q_t(n3087_t)
  );


  nnd2s3
  U1340
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n2278),
    .DIN2_t(n2278_t),
    .Q(n3086),
    .Q_t(n3086_t)
  );


  nnd2s3
  U1341
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n2267),
    .DIN2_t(n2267_t),
    .Q(n3085),
    .Q_t(n3085_t)
  );


  nnd2s3
  U1342
  (
    .DIN1(n6658),
    .DIN1_t(n6658_t),
    .DIN2(n3089),
    .DIN2_t(n3089_t),
    .Q(n3084),
    .Q_t(n3084_t)
  );


  nor2s3
  U1343
  (
    .DIN1(n5325),
    .DIN1_t(n5325_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6959),
    .Q_t(WX6959_t)
  );


  nor2s3
  U1344
  (
    .DIN1(n5326),
    .DIN1_t(n5326_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6957),
    .Q_t(WX6957_t)
  );


  nor2s3
  U1345
  (
    .DIN1(n5327),
    .DIN1_t(n5327_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6955),
    .Q_t(WX6955_t)
  );


  nor2s3
  U1346
  (
    .DIN1(n5328),
    .DIN1_t(n5328_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6953),
    .Q_t(WX6953_t)
  );


  nor2s3
  U1347
  (
    .DIN1(n5329),
    .DIN1_t(n5329_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6951),
    .Q_t(WX6951_t)
  );


  nor2s3
  U1348
  (
    .DIN1(n5330),
    .DIN1_t(n5330_t),
    .DIN2(n6713),
    .DIN2_t(n6713_t),
    .Q(WX6949),
    .Q_t(WX6949_t)
  );


  nnd4s2
  U1349
  (
    .DIN1(n3090),
    .DIN1_t(n3090_t),
    .DIN2(n3091),
    .DIN2_t(n3091_t),
    .DIN3(n3092),
    .DIN3_t(n3092_t),
    .DIN4(n3093),
    .DIN4_t(n3093_t),
    .Q(WX694),
    .Q_t(WX694_t)
  );


  nnd2s3
  U1350
  (
    .DIN1(n3094),
    .DIN1_t(n3094_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3093),
    .Q_t(n3093_t)
  );


  nnd2s3
  U1351
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n2279),
    .DIN2_t(n2279_t),
    .Q(n3092),
    .Q_t(n3092_t)
  );


  nnd2s3
  U1352
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n2266),
    .DIN2_t(n2266_t),
    .Q(n3091),
    .Q_t(n3091_t)
  );


  nnd2s3
  U1353
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3095),
    .DIN2_t(n3095_t),
    .Q(n3090),
    .Q_t(n3090_t)
  );


  nnd4s2
  U1354
  (
    .DIN1(n3096),
    .DIN1_t(n3096_t),
    .DIN2(n3097),
    .DIN2_t(n3097_t),
    .DIN3(n3098),
    .DIN3_t(n3098_t),
    .DIN4(n3099),
    .DIN4_t(n3099_t),
    .Q(WX692),
    .Q_t(WX692_t)
  );


  nnd2s3
  U1355
  (
    .DIN1(n3100),
    .DIN1_t(n3100_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3099),
    .Q_t(n3099_t)
  );


  nnd2s3
  U1356
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n2280),
    .DIN2_t(n2280_t),
    .Q(n3098),
    .Q_t(n3098_t)
  );


  nnd2s3
  U1357
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n2265),
    .DIN2_t(n2265_t),
    .Q(n3097),
    .Q_t(n3097_t)
  );


  nnd2s3
  U1358
  (
    .DIN1(n6658),
    .DIN1_t(n6658_t),
    .DIN2(n3101),
    .DIN2_t(n3101_t),
    .Q(n3096),
    .Q_t(n3096_t)
  );


  nnd4s2
  U1359
  (
    .DIN1(n3102),
    .DIN1_t(n3102_t),
    .DIN2(n3103),
    .DIN2_t(n3103_t),
    .DIN3(n3104),
    .DIN3_t(n3104_t),
    .DIN4(n3105),
    .DIN4_t(n3105_t),
    .Q(WX690),
    .Q_t(WX690_t)
  );


  nnd2s3
  U1360
  (
    .DIN1(n3106),
    .DIN1_t(n3106_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n3105),
    .Q_t(n3105_t)
  );


  nnd2s3
  U1361
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n2281),
    .DIN2_t(n2281_t),
    .Q(n3104),
    .Q_t(n3104_t)
  );


  nnd2s3
  U1362
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n2264),
    .DIN2_t(n2264_t),
    .Q(n3103),
    .Q_t(n3103_t)
  );


  nnd2s3
  U1363
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3107),
    .DIN2_t(n3107_t),
    .Q(n3102),
    .Q_t(n3102_t)
  );


  nnd4s2
  U1364
  (
    .DIN1(n3108),
    .DIN1_t(n3108_t),
    .DIN2(n3109),
    .DIN2_t(n3109_t),
    .DIN3(n3110),
    .DIN3_t(n3110_t),
    .DIN4(n3111),
    .DIN4_t(n3111_t),
    .Q(WX688),
    .Q_t(WX688_t)
  );


  nnd2s3
  U1365
  (
    .DIN1(n3112),
    .DIN1_t(n3112_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3111),
    .Q_t(n3111_t)
  );


  nnd2s3
  U1366
  (
    .DIN1(n6608),
    .DIN1_t(n6608_t),
    .DIN2(n2282),
    .DIN2_t(n2282_t),
    .Q(n3110),
    .Q_t(n3110_t)
  );


  nnd2s3
  U1367
  (
    .DIN1(n6577),
    .DIN1_t(n6577_t),
    .DIN2(n2263),
    .DIN2_t(n2263_t),
    .Q(n3109),
    .Q_t(n3109_t)
  );


  nnd2s3
  U1368
  (
    .DIN1(n6658),
    .DIN1_t(n6658_t),
    .DIN2(n3113),
    .DIN2_t(n3113_t),
    .Q(n3108),
    .Q_t(n3108_t)
  );


  nnd4s2
  U1369
  (
    .DIN1(n3114),
    .DIN1_t(n3114_t),
    .DIN2(n3115),
    .DIN2_t(n3115_t),
    .DIN3(n3116),
    .DIN3_t(n3116_t),
    .DIN4(n3117),
    .DIN4_t(n3117_t),
    .Q(WX686),
    .Q_t(WX686_t)
  );


  nnd2s3
  U1370
  (
    .DIN1(n3118),
    .DIN1_t(n3118_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3117),
    .Q_t(n3117_t)
  );


  nnd2s3
  U1371
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2283),
    .DIN2_t(n2283_t),
    .Q(n3116),
    .Q_t(n3116_t)
  );


  nnd2s3
  U1372
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2262),
    .DIN2_t(n2262_t),
    .Q(n3115),
    .Q_t(n3115_t)
  );


  nnd2s3
  U1373
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3119),
    .DIN2_t(n3119_t),
    .Q(n3114),
    .Q_t(n3114_t)
  );


  nnd4s2
  U1374
  (
    .DIN1(n3120),
    .DIN1_t(n3120_t),
    .DIN2(n3121),
    .DIN2_t(n3121_t),
    .DIN3(n3122),
    .DIN3_t(n3122_t),
    .DIN4(n3123),
    .DIN4_t(n3123_t),
    .Q(WX684),
    .Q_t(WX684_t)
  );


  nnd2s3
  U1375
  (
    .DIN1(n3124),
    .DIN1_t(n3124_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3123),
    .Q_t(n3123_t)
  );


  nnd2s3
  U1376
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2284),
    .DIN2_t(n2284_t),
    .Q(n3122),
    .Q_t(n3122_t)
  );


  nnd2s3
  U1377
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2261),
    .DIN2_t(n2261_t),
    .Q(n3121),
    .Q_t(n3121_t)
  );


  nnd2s3
  U1378
  (
    .DIN1(n6658),
    .DIN1_t(n6658_t),
    .DIN2(n3125),
    .DIN2_t(n3125_t),
    .Q(n3120),
    .Q_t(n3120_t)
  );


  nnd4s2
  U1379
  (
    .DIN1(n3126),
    .DIN1_t(n3126_t),
    .DIN2(n3127),
    .DIN2_t(n3127_t),
    .DIN3(n3128),
    .DIN3_t(n3128_t),
    .DIN4(n3129),
    .DIN4_t(n3129_t),
    .Q(WX682),
    .Q_t(WX682_t)
  );


  nnd2s3
  U1380
  (
    .DIN1(n3130),
    .DIN1_t(n3130_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3129),
    .Q_t(n3129_t)
  );


  nnd2s3
  U1381
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2285),
    .DIN2_t(n2285_t),
    .Q(n3128),
    .Q_t(n3128_t)
  );


  nnd2s3
  U1382
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2260),
    .DIN2_t(n2260_t),
    .Q(n3127),
    .Q_t(n3127_t)
  );


  nnd2s3
  U1383
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3131),
    .DIN2_t(n3131_t),
    .Q(n3126),
    .Q_t(n3126_t)
  );


  nnd4s2
  U1384
  (
    .DIN1(n3132),
    .DIN1_t(n3132_t),
    .DIN2(n3133),
    .DIN2_t(n3133_t),
    .DIN3(n3134),
    .DIN3_t(n3134_t),
    .DIN4(n3135),
    .DIN4_t(n3135_t),
    .Q(WX680),
    .Q_t(WX680_t)
  );


  nnd2s3
  U1385
  (
    .DIN1(n3136),
    .DIN1_t(n3136_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3135),
    .Q_t(n3135_t)
  );


  nnd2s3
  U1386
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2286),
    .DIN2_t(n2286_t),
    .Q(n3134),
    .Q_t(n3134_t)
  );


  nnd2s3
  U1387
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2259),
    .DIN2_t(n2259_t),
    .Q(n3133),
    .Q_t(n3133_t)
  );


  nnd2s3
  U1388
  (
    .DIN1(n6658),
    .DIN1_t(n6658_t),
    .DIN2(n3137),
    .DIN2_t(n3137_t),
    .Q(n3132),
    .Q_t(n3132_t)
  );


  nnd4s2
  U1389
  (
    .DIN1(n3138),
    .DIN1_t(n3138_t),
    .DIN2(n3139),
    .DIN2_t(n3139_t),
    .DIN3(n3140),
    .DIN3_t(n3140_t),
    .DIN4(n3141),
    .DIN4_t(n3141_t),
    .Q(WX678),
    .Q_t(WX678_t)
  );


  nnd2s3
  U1390
  (
    .DIN1(n3142),
    .DIN1_t(n3142_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3141),
    .Q_t(n3141_t)
  );


  nnd2s3
  U1391
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2287),
    .DIN2_t(n2287_t),
    .Q(n3140),
    .Q_t(n3140_t)
  );


  nnd2s3
  U1392
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2258),
    .DIN2_t(n2258_t),
    .Q(n3139),
    .Q_t(n3139_t)
  );


  nnd2s3
  U1393
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3143),
    .DIN2_t(n3143_t),
    .Q(n3138),
    .Q_t(n3138_t)
  );


  nnd4s2
  U1394
  (
    .DIN1(n3144),
    .DIN1_t(n3144_t),
    .DIN2(n3145),
    .DIN2_t(n3145_t),
    .DIN3(n3146),
    .DIN3_t(n3146_t),
    .DIN4(n3147),
    .DIN4_t(n3147_t),
    .Q(WX676),
    .Q_t(WX676_t)
  );


  nnd2s3
  U1395
  (
    .DIN1(n3148),
    .DIN1_t(n3148_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3147),
    .Q_t(n3147_t)
  );


  nnd2s3
  U1396
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2288),
    .DIN2_t(n2288_t),
    .Q(n3146),
    .Q_t(n3146_t)
  );


  nnd2s3
  U1397
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2257),
    .DIN2_t(n2257_t),
    .Q(n3145),
    .Q_t(n3145_t)
  );


  nnd2s3
  U1398
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3149),
    .DIN2_t(n3149_t),
    .Q(n3144),
    .Q_t(n3144_t)
  );


  nnd4s2
  U1399
  (
    .DIN1(n3150),
    .DIN1_t(n3150_t),
    .DIN2(n3151),
    .DIN2_t(n3151_t),
    .DIN3(n3152),
    .DIN3_t(n3152_t),
    .DIN4(n3153),
    .DIN4_t(n3153_t),
    .Q(WX674),
    .Q_t(WX674_t)
  );


  nnd2s3
  U1400
  (
    .DIN1(n3154),
    .DIN1_t(n3154_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3153),
    .Q_t(n3153_t)
  );


  nnd2s3
  U1401
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2289),
    .DIN2_t(n2289_t),
    .Q(n3152),
    .Q_t(n3152_t)
  );


  nnd2s3
  U1402
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2256),
    .DIN2_t(n2256_t),
    .Q(n3151),
    .Q_t(n3151_t)
  );


  nnd2s3
  U1403
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3155),
    .DIN2_t(n3155_t),
    .Q(n3150),
    .Q_t(n3150_t)
  );


  nnd4s2
  U1404
  (
    .DIN1(n3156),
    .DIN1_t(n3156_t),
    .DIN2(n3157),
    .DIN2_t(n3157_t),
    .DIN3(n3158),
    .DIN3_t(n3158_t),
    .DIN4(n3159),
    .DIN4_t(n3159_t),
    .Q(WX672),
    .Q_t(WX672_t)
  );


  nnd2s3
  U1405
  (
    .DIN1(n3160),
    .DIN1_t(n3160_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3159),
    .Q_t(n3159_t)
  );


  nnd2s3
  U1406
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2290),
    .DIN2_t(n2290_t),
    .Q(n3158),
    .Q_t(n3158_t)
  );


  nnd2s3
  U1407
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2255),
    .DIN2_t(n2255_t),
    .Q(n3157),
    .Q_t(n3157_t)
  );


  nnd2s3
  U1408
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3161),
    .DIN2_t(n3161_t),
    .Q(n3156),
    .Q_t(n3156_t)
  );


  nnd4s2
  U1409
  (
    .DIN1(n3162),
    .DIN1_t(n3162_t),
    .DIN2(n3163),
    .DIN2_t(n3163_t),
    .DIN3(n3164),
    .DIN3_t(n3164_t),
    .DIN4(n3165),
    .DIN4_t(n3165_t),
    .Q(WX670),
    .Q_t(WX670_t)
  );


  nnd2s3
  U1410
  (
    .DIN1(n3166),
    .DIN1_t(n3166_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3165),
    .Q_t(n3165_t)
  );


  nnd2s3
  U1411
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2291),
    .DIN2_t(n2291_t),
    .Q(n3164),
    .Q_t(n3164_t)
  );


  nnd2s3
  U1412
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2254),
    .DIN2_t(n2254_t),
    .Q(n3163),
    .Q_t(n3163_t)
  );


  nnd2s3
  U1413
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3167),
    .DIN2_t(n3167_t),
    .Q(n3162),
    .Q_t(n3162_t)
  );


  nnd4s2
  U1414
  (
    .DIN1(n3168),
    .DIN1_t(n3168_t),
    .DIN2(n3169),
    .DIN2_t(n3169_t),
    .DIN3(n3170),
    .DIN3_t(n3170_t),
    .DIN4(n3171),
    .DIN4_t(n3171_t),
    .Q(WX668),
    .Q_t(WX668_t)
  );


  nnd2s3
  U1415
  (
    .DIN1(n3172),
    .DIN1_t(n3172_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3171),
    .Q_t(n3171_t)
  );


  nnd2s3
  U1416
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2292),
    .DIN2_t(n2292_t),
    .Q(n3170),
    .Q_t(n3170_t)
  );


  nnd2s3
  U1417
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2253),
    .DIN2_t(n2253_t),
    .Q(n3169),
    .Q_t(n3169_t)
  );


  nnd2s3
  U1418
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3173),
    .DIN2_t(n3173_t),
    .Q(n3168),
    .Q_t(n3168_t)
  );


  nnd4s2
  U1419
  (
    .DIN1(n3174),
    .DIN1_t(n3174_t),
    .DIN2(n3175),
    .DIN2_t(n3175_t),
    .DIN3(n3176),
    .DIN3_t(n3176_t),
    .DIN4(n3177),
    .DIN4_t(n3177_t),
    .Q(WX666),
    .Q_t(WX666_t)
  );


  nnd2s3
  U1420
  (
    .DIN1(n3178),
    .DIN1_t(n3178_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3177),
    .Q_t(n3177_t)
  );


  nnd2s3
  U1421
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2293),
    .DIN2_t(n2293_t),
    .Q(n3176),
    .Q_t(n3176_t)
  );


  nnd2s3
  U1422
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2252),
    .DIN2_t(n2252_t),
    .Q(n3175),
    .Q_t(n3175_t)
  );


  nnd2s3
  U1423
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3179),
    .DIN2_t(n3179_t),
    .Q(n3174),
    .Q_t(n3174_t)
  );


  nnd4s2
  U1424
  (
    .DIN1(n3180),
    .DIN1_t(n3180_t),
    .DIN2(n3181),
    .DIN2_t(n3181_t),
    .DIN3(n3182),
    .DIN3_t(n3182_t),
    .DIN4(n3183),
    .DIN4_t(n3183_t),
    .Q(WX664),
    .Q_t(WX664_t)
  );


  nnd2s3
  U1425
  (
    .DIN1(n3184),
    .DIN1_t(n3184_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3183),
    .Q_t(n3183_t)
  );


  nnd2s3
  U1426
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2294),
    .DIN2_t(n2294_t),
    .Q(n3182),
    .Q_t(n3182_t)
  );


  nnd2s3
  U1427
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2251),
    .DIN2_t(n2251_t),
    .Q(n3181),
    .Q_t(n3181_t)
  );


  nnd2s3
  U1428
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3185),
    .DIN2_t(n3185_t),
    .Q(n3180),
    .Q_t(n3180_t)
  );


  nnd4s2
  U1429
  (
    .DIN1(n3186),
    .DIN1_t(n3186_t),
    .DIN2(n3187),
    .DIN2_t(n3187_t),
    .DIN3(n3188),
    .DIN3_t(n3188_t),
    .DIN4(n3189),
    .DIN4_t(n3189_t),
    .Q(WX662),
    .Q_t(WX662_t)
  );


  nnd2s3
  U1430
  (
    .DIN1(n3190),
    .DIN1_t(n3190_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3189),
    .Q_t(n3189_t)
  );


  nnd2s3
  U1431
  (
    .DIN1(n6607),
    .DIN1_t(n6607_t),
    .DIN2(n2295),
    .DIN2_t(n2295_t),
    .Q(n3188),
    .Q_t(n3188_t)
  );


  nnd2s3
  U1432
  (
    .DIN1(n6576),
    .DIN1_t(n6576_t),
    .DIN2(n2250),
    .DIN2_t(n2250_t),
    .Q(n3187),
    .Q_t(n3187_t)
  );


  nnd2s3
  U1433
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3191),
    .DIN2_t(n3191_t),
    .Q(n3186),
    .Q_t(n3186_t)
  );


  nnd4s2
  U1434
  (
    .DIN1(n3192),
    .DIN1_t(n3192_t),
    .DIN2(n3193),
    .DIN2_t(n3193_t),
    .DIN3(n3194),
    .DIN3_t(n3194_t),
    .DIN4(n3195),
    .DIN4_t(n3195_t),
    .Q(WX660),
    .Q_t(WX660_t)
  );


  nnd2s3
  U1435
  (
    .DIN1(n3196),
    .DIN1_t(n3196_t),
    .DIN2(n6627),
    .DIN2_t(n6627_t),
    .Q(n3195),
    .Q_t(n3195_t)
  );


  nnd2s3
  U1436
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2296),
    .DIN2_t(n2296_t),
    .Q(n3194),
    .Q_t(n3194_t)
  );


  nnd2s3
  U1437
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2249),
    .DIN2_t(n2249_t),
    .Q(n3193),
    .Q_t(n3193_t)
  );


  nnd2s3
  U1438
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3197),
    .DIN2_t(n3197_t),
    .Q(n3192),
    .Q_t(n3192_t)
  );


  nnd4s2
  U1439
  (
    .DIN1(n3198),
    .DIN1_t(n3198_t),
    .DIN2(n3199),
    .DIN2_t(n3199_t),
    .DIN3(n3200),
    .DIN3_t(n3200_t),
    .DIN4(n3201),
    .DIN4_t(n3201_t),
    .Q(WX658),
    .Q_t(WX658_t)
  );


  nnd2s3
  U1440
  (
    .DIN1(n3202),
    .DIN1_t(n3202_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3201),
    .Q_t(n3201_t)
  );


  nnd2s3
  U1441
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2297),
    .DIN2_t(n2297_t),
    .Q(n3200),
    .Q_t(n3200_t)
  );


  nnd2s3
  U1442
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2248),
    .DIN2_t(n2248_t),
    .Q(n3199),
    .Q_t(n3199_t)
  );


  nnd2s3
  U1443
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3203),
    .DIN2_t(n3203_t),
    .Q(n3198),
    .Q_t(n3198_t)
  );


  nnd4s2
  U1444
  (
    .DIN1(n3204),
    .DIN1_t(n3204_t),
    .DIN2(n3333),
    .DIN2_t(n3333_t),
    .DIN3(n3334),
    .DIN3_t(n3334_t),
    .DIN4(n3335),
    .DIN4_t(n3335_t),
    .Q(WX656),
    .Q_t(WX656_t)
  );


  nnd2s3
  U1445
  (
    .DIN1(n3336),
    .DIN1_t(n3336_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3335),
    .Q_t(n3335_t)
  );


  nnd2s3
  U1446
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2298),
    .DIN2_t(n2298_t),
    .Q(n3334),
    .Q_t(n3334_t)
  );


  nnd2s3
  U1447
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2247),
    .DIN2_t(n2247_t),
    .Q(n3333),
    .Q_t(n3333_t)
  );


  nnd2s3
  U1448
  (
    .DIN1(n6657),
    .DIN1_t(n6657_t),
    .DIN2(n3337),
    .DIN2_t(n3337_t),
    .Q(n3204),
    .Q_t(n3204_t)
  );


  nnd4s2
  U1449
  (
    .DIN1(n3338),
    .DIN1_t(n3338_t),
    .DIN2(n3339),
    .DIN2_t(n3339_t),
    .DIN3(n3340),
    .DIN3_t(n3340_t),
    .DIN4(n3341),
    .DIN4_t(n3341_t),
    .Q(WX654),
    .Q_t(WX654_t)
  );


  nnd2s3
  U1450
  (
    .DIN1(n3342),
    .DIN1_t(n3342_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3341),
    .Q_t(n3341_t)
  );


  nnd2s3
  U1451
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2299),
    .DIN2_t(n2299_t),
    .Q(n3340),
    .Q_t(n3340_t)
  );


  nnd2s3
  U1452
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2246),
    .DIN2_t(n2246_t),
    .Q(n3339),
    .Q_t(n3339_t)
  );


  nnd2s3
  U1453
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3343),
    .DIN2_t(n3343_t),
    .Q(n3338),
    .Q_t(n3338_t)
  );


  nnd4s2
  U1454
  (
    .DIN1(n3344),
    .DIN1_t(n3344_t),
    .DIN2(n3345),
    .DIN2_t(n3345_t),
    .DIN3(n3346),
    .DIN3_t(n3346_t),
    .DIN4(n3347),
    .DIN4_t(n3347_t),
    .Q(WX652),
    .Q_t(WX652_t)
  );


  nnd2s3
  U1455
  (
    .DIN1(n3348),
    .DIN1_t(n3348_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3347),
    .Q_t(n3347_t)
  );


  nnd2s3
  U1456
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2300),
    .DIN2_t(n2300_t),
    .Q(n3346),
    .Q_t(n3346_t)
  );


  nnd2s3
  U1457
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2245),
    .DIN2_t(n2245_t),
    .Q(n3345),
    .Q_t(n3345_t)
  );


  nnd2s3
  U1458
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3349),
    .DIN2_t(n3349_t),
    .Q(n3344),
    .Q_t(n3344_t)
  );


  nnd4s2
  U1459
  (
    .DIN1(n3350),
    .DIN1_t(n3350_t),
    .DIN2(n3351),
    .DIN2_t(n3351_t),
    .DIN3(n3352),
    .DIN3_t(n3352_t),
    .DIN4(n3353),
    .DIN4_t(n3353_t),
    .Q(WX650),
    .Q_t(WX650_t)
  );


  nnd2s3
  U1460
  (
    .DIN1(n3354),
    .DIN1_t(n3354_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3353),
    .Q_t(n3353_t)
  );


  nnd2s3
  U1461
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2301),
    .DIN2_t(n2301_t),
    .Q(n3352),
    .Q_t(n3352_t)
  );


  nnd2s3
  U1462
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2244),
    .DIN2_t(n2244_t),
    .Q(n3351),
    .Q_t(n3351_t)
  );


  nnd2s3
  U1463
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3355),
    .DIN2_t(n3355_t),
    .Q(n3350),
    .Q_t(n3350_t)
  );


  nor2s3
  U1464
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n3356),
    .DIN2_t(n3356_t),
    .Q(WX6498),
    .Q_t(WX6498_t)
  );


  xor2s3
  U1465
  (
    .DIN1(n5469),
    .DIN1_t(n5469_t),
    .DIN2(n5649),
    .DIN2_t(n5649_t),
    .Q(n3356),
    .Q_t(n3356_t)
  );


  nor2s3
  U1466
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n3357),
    .DIN2_t(n3357_t),
    .Q(WX6496),
    .Q_t(WX6496_t)
  );


  xor2s3
  U1467
  (
    .DIN1(n5464),
    .DIN1_t(n5464_t),
    .DIN2(n5644),
    .DIN2_t(n5644_t),
    .Q(n3357),
    .Q_t(n3357_t)
  );


  nor2s3
  U1468
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n3358),
    .DIN2_t(n3358_t),
    .Q(WX6494),
    .Q_t(WX6494_t)
  );


  xor2s3
  U1469
  (
    .DIN1(n5459),
    .DIN1_t(n5459_t),
    .DIN2(n5639),
    .DIN2_t(n5639_t),
    .Q(n3358),
    .Q_t(n3358_t)
  );


  nor2s3
  U1470
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n3359),
    .DIN2_t(n3359_t),
    .Q(WX6492),
    .Q_t(WX6492_t)
  );


  xor2s3
  U1471
  (
    .DIN1(n5454),
    .DIN1_t(n5454_t),
    .DIN2(n5634),
    .DIN2_t(n5634_t),
    .Q(n3359),
    .Q_t(n3359_t)
  );


  nor2s3
  U1472
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n3360),
    .DIN2_t(n3360_t),
    .Q(WX6490),
    .Q_t(WX6490_t)
  );


  xor2s3
  U1473
  (
    .DIN1(n5449),
    .DIN1_t(n5449_t),
    .DIN2(n5629),
    .DIN2_t(n5629_t),
    .Q(n3360),
    .Q_t(n3360_t)
  );


  nor2s3
  U1474
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n3361),
    .DIN2_t(n3361_t),
    .Q(WX6488),
    .Q_t(WX6488_t)
  );


  xor2s3
  U1475
  (
    .DIN1(n5444),
    .DIN1_t(n5444_t),
    .DIN2(n5624),
    .DIN2_t(n5624_t),
    .Q(n3361),
    .Q_t(n3361_t)
  );


  nor2s3
  U1476
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n3362),
    .DIN2_t(n3362_t),
    .Q(WX6486),
    .Q_t(WX6486_t)
  );


  xor2s3
  U1477
  (
    .DIN1(n5439),
    .DIN1_t(n5439_t),
    .DIN2(n5619),
    .DIN2_t(n5619_t),
    .Q(n3362),
    .Q_t(n3362_t)
  );


  nor2s3
  U1478
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n3363),
    .DIN2_t(n3363_t),
    .Q(WX6484),
    .Q_t(WX6484_t)
  );


  xor2s3
  U1479
  (
    .DIN1(n5434),
    .DIN1_t(n5434_t),
    .DIN2(n5614),
    .DIN2_t(n5614_t),
    .Q(n3363),
    .Q_t(n3363_t)
  );


  nor2s3
  U1480
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n3364),
    .DIN2_t(n3364_t),
    .Q(WX6482),
    .Q_t(WX6482_t)
  );


  xor2s3
  U1481
  (
    .DIN1(n5429),
    .DIN1_t(n5429_t),
    .DIN2(n5609),
    .DIN2_t(n5609_t),
    .Q(n3364),
    .Q_t(n3364_t)
  );


  nor2s3
  U1482
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n3365),
    .DIN2_t(n3365_t),
    .Q(WX6480),
    .Q_t(WX6480_t)
  );


  xor2s3
  U1483
  (
    .DIN1(n5424),
    .DIN1_t(n5424_t),
    .DIN2(n5604),
    .DIN2_t(n5604_t),
    .Q(n3365),
    .Q_t(n3365_t)
  );


  nnd4s2
  U1484
  (
    .DIN1(n3366),
    .DIN1_t(n3366_t),
    .DIN2(n3367),
    .DIN2_t(n3367_t),
    .DIN3(n3368),
    .DIN3_t(n3368_t),
    .DIN4(n3369),
    .DIN4_t(n3369_t),
    .Q(WX648),
    .Q_t(WX648_t)
  );


  nnd2s3
  U1485
  (
    .DIN1(n3370),
    .DIN1_t(n3370_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3369),
    .Q_t(n3369_t)
  );


  nnd2s3
  U1486
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2302),
    .DIN2_t(n2302_t),
    .Q(n3368),
    .Q_t(n3368_t)
  );


  nnd2s3
  U1487
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2243),
    .DIN2_t(n2243_t),
    .Q(n3367),
    .Q_t(n3367_t)
  );


  nnd2s3
  U1488
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3371),
    .DIN2_t(n3371_t),
    .Q(n3366),
    .Q_t(n3366_t)
  );


  nor2s3
  U1489
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3372),
    .DIN2_t(n3372_t),
    .Q(WX6478),
    .Q_t(WX6478_t)
  );


  xor2s3
  U1490
  (
    .DIN1(n5419),
    .DIN1_t(n5419_t),
    .DIN2(n5599),
    .DIN2_t(n5599_t),
    .Q(n3372),
    .Q_t(n3372_t)
  );


  nor2s3
  U1491
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3373),
    .DIN2_t(n3373_t),
    .Q(WX6476),
    .Q_t(WX6476_t)
  );


  xor2s3
  U1492
  (
    .DIN1(n5414),
    .DIN1_t(n5414_t),
    .DIN2(n5594),
    .DIN2_t(n5594_t),
    .Q(n3373),
    .Q_t(n3373_t)
  );


  nor2s3
  U1493
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3374),
    .DIN2_t(n3374_t),
    .Q(WX6474),
    .Q_t(WX6474_t)
  );


  xor2s3
  U1494
  (
    .DIN1(n5409),
    .DIN1_t(n5409_t),
    .DIN2(n5589),
    .DIN2_t(n5589_t),
    .Q(n3374),
    .Q_t(n3374_t)
  );


  nor2s3
  U1495
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3375),
    .DIN2_t(n3375_t),
    .Q(WX6472),
    .Q_t(WX6472_t)
  );


  xor2s3
  U1496
  (
    .DIN1(n5404),
    .DIN1_t(n5404_t),
    .DIN2(n5584),
    .DIN2_t(n5584_t),
    .Q(n3375),
    .Q_t(n3375_t)
  );


  nor2s3
  U1497
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3376),
    .DIN2_t(n3376_t),
    .Q(WX6470),
    .Q_t(WX6470_t)
  );


  xor2s3
  U1498
  (
    .DIN1(n5399),
    .DIN1_t(n5399_t),
    .DIN2(n5579),
    .DIN2_t(n5579_t),
    .Q(n3376),
    .Q_t(n3376_t)
  );


  nor2s3
  U1499
  (
    .DIN1(n3377),
    .DIN1_t(n3377_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX6468),
    .Q_t(WX6468_t)
  );


  xnr2s3
  U1500
  (
    .DIN1(n5574),
    .DIN1_t(n5574_t),
    .DIN2(n3378),
    .DIN2_t(n3378_t),
    .Q(n3377),
    .Q_t(n3377_t)
  );


  xor2s3
  U1501
  (
    .DIN1(n5394),
    .DIN1_t(n5394_t),
    .DIN2(n5474),
    .DIN2_t(n5474_t),
    .Q(n3378),
    .Q_t(n3378_t)
  );


  nor2s3
  U1502
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3379),
    .DIN2_t(n3379_t),
    .Q(WX6466),
    .Q_t(WX6466_t)
  );


  xor2s3
  U1503
  (
    .DIN1(n5390),
    .DIN1_t(n5390_t),
    .DIN2(n3268),
    .DIN2_t(n3268_t),
    .Q(n3379),
    .Q_t(n3379_t)
  );


  nor2s3
  U1504
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3380),
    .DIN2_t(n3380_t),
    .Q(WX6464),
    .Q_t(WX6464_t)
  );


  xor2s3
  U1505
  (
    .DIN1(n5386),
    .DIN1_t(n5386_t),
    .DIN2(n3267),
    .DIN2_t(n3267_t),
    .Q(n3380),
    .Q_t(n3380_t)
  );


  nor2s3
  U1506
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3381),
    .DIN2_t(n3381_t),
    .Q(WX6462),
    .Q_t(WX6462_t)
  );


  xor2s3
  U1507
  (
    .DIN1(n5382),
    .DIN1_t(n5382_t),
    .DIN2(n3266),
    .DIN2_t(n3266_t),
    .Q(n3381),
    .Q_t(n3381_t)
  );


  nor2s3
  U1508
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3382),
    .DIN2_t(n3382_t),
    .Q(WX6460),
    .Q_t(WX6460_t)
  );


  xor2s3
  U1509
  (
    .DIN1(n5378),
    .DIN1_t(n5378_t),
    .DIN2(n3265),
    .DIN2_t(n3265_t),
    .Q(n3382),
    .Q_t(n3382_t)
  );


  nnd4s2
  U1510
  (
    .DIN1(n3383),
    .DIN1_t(n3383_t),
    .DIN2(n3384),
    .DIN2_t(n3384_t),
    .DIN3(n3385),
    .DIN3_t(n3385_t),
    .DIN4(n3386),
    .DIN4_t(n3386_t),
    .Q(WX646),
    .Q_t(WX646_t)
  );


  nnd2s3
  U1511
  (
    .DIN1(n3387),
    .DIN1_t(n3387_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3386),
    .Q_t(n3386_t)
  );


  nnd2s3
  U1512
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2303),
    .DIN2_t(n2303_t),
    .Q(n3385),
    .Q_t(n3385_t)
  );


  nnd2s3
  U1513
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2242),
    .DIN2_t(n2242_t),
    .Q(n3384),
    .Q_t(n3384_t)
  );


  nnd2s3
  U1514
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3388),
    .DIN2_t(n3388_t),
    .Q(n3383),
    .Q_t(n3383_t)
  );


  nor2s3
  U1515
  (
    .DIN1(n3389),
    .DIN1_t(n3389_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX6458),
    .Q_t(WX6458_t)
  );


  xnr2s3
  U1516
  (
    .DIN1(n3264),
    .DIN1_t(n3264_t),
    .DIN2(n3390),
    .DIN2_t(n3390_t),
    .Q(n3389),
    .Q_t(n3389_t)
  );


  xor2s3
  U1517
  (
    .DIN1(n5374),
    .DIN1_t(n5374_t),
    .DIN2(n5474),
    .DIN2_t(n5474_t),
    .Q(n3390),
    .Q_t(n3390_t)
  );


  nor2s3
  U1518
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3391),
    .DIN2_t(n3391_t),
    .Q(WX6456),
    .Q_t(WX6456_t)
  );


  xor2s3
  U1519
  (
    .DIN1(n5370),
    .DIN1_t(n5370_t),
    .DIN2(n3263),
    .DIN2_t(n3263_t),
    .Q(n3391),
    .Q_t(n3391_t)
  );


  nor2s3
  U1520
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3392),
    .DIN2_t(n3392_t),
    .Q(WX6454),
    .Q_t(WX6454_t)
  );


  xor2s3
  U1521
  (
    .DIN1(n5366),
    .DIN1_t(n5366_t),
    .DIN2(n3262),
    .DIN2_t(n3262_t),
    .Q(n3392),
    .Q_t(n3392_t)
  );


  nor2s3
  U1522
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3393),
    .DIN2_t(n3393_t),
    .Q(WX6452),
    .Q_t(WX6452_t)
  );


  xor2s3
  U1523
  (
    .DIN1(n5362),
    .DIN1_t(n5362_t),
    .DIN2(n3261),
    .DIN2_t(n3261_t),
    .Q(n3393),
    .Q_t(n3393_t)
  );


  nor2s3
  U1524
  (
    .DIN1(n6799),
    .DIN1_t(n6799_t),
    .DIN2(n3394),
    .DIN2_t(n3394_t),
    .Q(WX6450),
    .Q_t(WX6450_t)
  );


  xor2s3
  U1525
  (
    .DIN1(n5358),
    .DIN1_t(n5358_t),
    .DIN2(n3260),
    .DIN2_t(n3260_t),
    .Q(n3394),
    .Q_t(n3394_t)
  );


  nor2s3
  U1526
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n3395),
    .DIN2_t(n3395_t),
    .Q(WX6448),
    .Q_t(WX6448_t)
  );


  xor2s3
  U1527
  (
    .DIN1(n5354),
    .DIN1_t(n5354_t),
    .DIN2(n3259),
    .DIN2_t(n3259_t),
    .Q(n3395),
    .Q_t(n3395_t)
  );


  nor2s3
  U1528
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n3396),
    .DIN2_t(n3396_t),
    .Q(WX6446),
    .Q_t(WX6446_t)
  );


  xor2s3
  U1529
  (
    .DIN1(n5350),
    .DIN1_t(n5350_t),
    .DIN2(n3258),
    .DIN2_t(n3258_t),
    .Q(n3396),
    .Q_t(n3396_t)
  );


  nor2s3
  U1530
  (
    .DIN1(n3397),
    .DIN1_t(n3397_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX6444),
    .Q_t(WX6444_t)
  );


  xnr2s3
  U1531
  (
    .DIN1(n3257),
    .DIN1_t(n3257_t),
    .DIN2(n3398),
    .DIN2_t(n3398_t),
    .Q(n3397),
    .Q_t(n3397_t)
  );


  xor2s3
  U1532
  (
    .DIN1(n5346),
    .DIN1_t(n5346_t),
    .DIN2(n5474),
    .DIN2_t(n5474_t),
    .Q(n3398),
    .Q_t(n3398_t)
  );


  nor2s3
  U1533
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n3399),
    .DIN2_t(n3399_t),
    .Q(WX6442),
    .Q_t(WX6442_t)
  );


  xor2s3
  U1534
  (
    .DIN1(n5342),
    .DIN1_t(n5342_t),
    .DIN2(n3256),
    .DIN2_t(n3256_t),
    .Q(n3399),
    .Q_t(n3399_t)
  );


  nor2s3
  U1535
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n3400),
    .DIN2_t(n3400_t),
    .Q(WX6440),
    .Q_t(WX6440_t)
  );


  xor2s3
  U1536
  (
    .DIN1(n5338),
    .DIN1_t(n5338_t),
    .DIN2(n3255),
    .DIN2_t(n3255_t),
    .Q(n3400),
    .Q_t(n3400_t)
  );


  nnd4s2
  U1537
  (
    .DIN1(n3401),
    .DIN1_t(n3401_t),
    .DIN2(n3402),
    .DIN2_t(n3402_t),
    .DIN3(n3403),
    .DIN3_t(n3403_t),
    .DIN4(n3404),
    .DIN4_t(n3404_t),
    .Q(WX644),
    .Q_t(WX644_t)
  );


  nnd2s3
  U1538
  (
    .DIN1(n3405),
    .DIN1_t(n3405_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3404),
    .Q_t(n3404_t)
  );


  nnd2s3
  U1539
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2304),
    .DIN2_t(n2304_t),
    .Q(n3403),
    .Q_t(n3403_t)
  );


  nnd2s3
  U1540
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2241),
    .DIN2_t(n2241_t),
    .Q(n3402),
    .Q_t(n3402_t)
  );


  nnd2s3
  U1541
  (
    .DIN1(n6656),
    .DIN1_t(n6656_t),
    .DIN2(n3406),
    .DIN2_t(n3406_t),
    .Q(n3401),
    .Q_t(n3401_t)
  );


  nor2s3
  U1542
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n3407),
    .DIN2_t(n3407_t),
    .Q(WX6438),
    .Q_t(WX6438_t)
  );


  xor2s3
  U1543
  (
    .DIN1(n5334),
    .DIN1_t(n5334_t),
    .DIN2(n3254),
    .DIN2_t(n3254_t),
    .Q(n3407),
    .Q_t(n3407_t)
  );


  nor2s3
  U1544
  (
    .DIN1(n6800),
    .DIN1_t(n6800_t),
    .DIN2(n3408),
    .DIN2_t(n3408_t),
    .Q(WX6436),
    .Q_t(WX6436_t)
  );


  xor2s3
  U1545
  (
    .DIN1(n5474),
    .DIN1_t(n5474_t),
    .DIN2(n3253),
    .DIN2_t(n3253_t),
    .Q(n3408),
    .Q_t(n3408_t)
  );


  nor2s3
  U1546
  (
    .DIN1(n5509),
    .DIN1_t(n5509_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX6070),
    .Q_t(WX6070_t)
  );


  nor2s3
  U1547
  (
    .DIN1(n5513),
    .DIN1_t(n5513_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX6068),
    .Q_t(WX6068_t)
  );


  nor2s3
  U1548
  (
    .DIN1(n5517),
    .DIN1_t(n5517_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX6066),
    .Q_t(WX6066_t)
  );


  nor2s3
  U1549
  (
    .DIN1(n5521),
    .DIN1_t(n5521_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX6064),
    .Q_t(WX6064_t)
  );


  nor2s3
  U1550
  (
    .DIN1(n5525),
    .DIN1_t(n5525_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX6062),
    .Q_t(WX6062_t)
  );


  nor2s3
  U1551
  (
    .DIN1(n5529),
    .DIN1_t(n5529_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX6060),
    .Q_t(WX6060_t)
  );


  nor2s3
  U1552
  (
    .DIN1(n5533),
    .DIN1_t(n5533_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX6058),
    .Q_t(WX6058_t)
  );


  nor2s3
  U1553
  (
    .DIN1(n5537),
    .DIN1_t(n5537_t),
    .DIN2(n6712),
    .DIN2_t(n6712_t),
    .Q(WX6056),
    .Q_t(WX6056_t)
  );


  nor2s3
  U1554
  (
    .DIN1(n5541),
    .DIN1_t(n5541_t),
    .DIN2(n6717),
    .DIN2_t(n6717_t),
    .Q(WX6054),
    .Q_t(WX6054_t)
  );


  nor2s3
  U1555
  (
    .DIN1(n5545),
    .DIN1_t(n5545_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX6052),
    .Q_t(WX6052_t)
  );


  nor2s3
  U1556
  (
    .DIN1(n5549),
    .DIN1_t(n5549_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6050),
    .Q_t(WX6050_t)
  );


  nor2s3
  U1557
  (
    .DIN1(n5553),
    .DIN1_t(n5553_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6048),
    .Q_t(WX6048_t)
  );


  nor2s3
  U1558
  (
    .DIN1(n5557),
    .DIN1_t(n5557_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6046),
    .Q_t(WX6046_t)
  );


  nor2s3
  U1559
  (
    .DIN1(n5561),
    .DIN1_t(n5561_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6044),
    .Q_t(WX6044_t)
  );


  nor2s3
  U1560
  (
    .DIN1(n5565),
    .DIN1_t(n5565_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6042),
    .Q_t(WX6042_t)
  );


  nor2s3
  U1561
  (
    .DIN1(n5569),
    .DIN1_t(n5569_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6040),
    .Q_t(WX6040_t)
  );


  nor2s3
  U1562
  (
    .DIN1(n5573),
    .DIN1_t(n5573_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6038),
    .Q_t(WX6038_t)
  );


  nor2s3
  U1563
  (
    .DIN1(n5578),
    .DIN1_t(n5578_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6036),
    .Q_t(WX6036_t)
  );


  nor2s3
  U1564
  (
    .DIN1(n5583),
    .DIN1_t(n5583_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6034),
    .Q_t(WX6034_t)
  );


  nor2s3
  U1565
  (
    .DIN1(n5588),
    .DIN1_t(n5588_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6032),
    .Q_t(WX6032_t)
  );


  nor2s3
  U1566
  (
    .DIN1(n5593),
    .DIN1_t(n5593_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6030),
    .Q_t(WX6030_t)
  );


  nor2s3
  U1567
  (
    .DIN1(n5598),
    .DIN1_t(n5598_t),
    .DIN2(n6733),
    .DIN2_t(n6733_t),
    .Q(WX6028),
    .Q_t(WX6028_t)
  );


  nor2s3
  U1568
  (
    .DIN1(n5603),
    .DIN1_t(n5603_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6026),
    .Q_t(WX6026_t)
  );


  nor2s3
  U1569
  (
    .DIN1(n5608),
    .DIN1_t(n5608_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6024),
    .Q_t(WX6024_t)
  );


  nor2s3
  U1570
  (
    .DIN1(n5613),
    .DIN1_t(n5613_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6022),
    .Q_t(WX6022_t)
  );


  nor2s3
  U1571
  (
    .DIN1(n5618),
    .DIN1_t(n5618_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6020),
    .Q_t(WX6020_t)
  );


  nor2s3
  U1572
  (
    .DIN1(n5623),
    .DIN1_t(n5623_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6018),
    .Q_t(WX6018_t)
  );


  nor2s3
  U1573
  (
    .DIN1(n5628),
    .DIN1_t(n5628_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6016),
    .Q_t(WX6016_t)
  );


  nor2s3
  U1574
  (
    .DIN1(n5633),
    .DIN1_t(n5633_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6014),
    .Q_t(WX6014_t)
  );


  nor2s3
  U1575
  (
    .DIN1(n5638),
    .DIN1_t(n5638_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6012),
    .Q_t(WX6012_t)
  );


  nor2s3
  U1576
  (
    .DIN1(n5643),
    .DIN1_t(n5643_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6010),
    .Q_t(WX6010_t)
  );


  nor2s3
  U1577
  (
    .DIN1(n5648),
    .DIN1_t(n5648_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6008),
    .Q_t(WX6008_t)
  );


  nor2s3
  U1578
  (
    .DIN1(n5508),
    .DIN1_t(n5508_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6006),
    .Q_t(WX6006_t)
  );


  nor2s3
  U1579
  (
    .DIN1(n5512),
    .DIN1_t(n5512_t),
    .DIN2(n6732),
    .DIN2_t(n6732_t),
    .Q(WX6004),
    .Q_t(WX6004_t)
  );


  nor2s3
  U1580
  (
    .DIN1(n5516),
    .DIN1_t(n5516_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX6002),
    .Q_t(WX6002_t)
  );


  nor2s3
  U1581
  (
    .DIN1(n5520),
    .DIN1_t(n5520_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX6000),
    .Q_t(WX6000_t)
  );


  nor2s3
  U1582
  (
    .DIN1(n5524),
    .DIN1_t(n5524_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX5998),
    .Q_t(WX5998_t)
  );


  nor2s3
  U1583
  (
    .DIN1(n5528),
    .DIN1_t(n5528_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX5996),
    .Q_t(WX5996_t)
  );


  nor2s3
  U1584
  (
    .DIN1(n5532),
    .DIN1_t(n5532_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX5994),
    .Q_t(WX5994_t)
  );


  nor2s3
  U1585
  (
    .DIN1(n5536),
    .DIN1_t(n5536_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX5992),
    .Q_t(WX5992_t)
  );


  nor2s3
  U1586
  (
    .DIN1(n5540),
    .DIN1_t(n5540_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX5990),
    .Q_t(WX5990_t)
  );


  nor2s3
  U1587
  (
    .DIN1(n5544),
    .DIN1_t(n5544_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX5988),
    .Q_t(WX5988_t)
  );


  nor2s3
  U1588
  (
    .DIN1(n5548),
    .DIN1_t(n5548_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX5986),
    .Q_t(WX5986_t)
  );


  nor2s3
  U1589
  (
    .DIN1(n5552),
    .DIN1_t(n5552_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX5984),
    .Q_t(WX5984_t)
  );


  nor2s3
  U1590
  (
    .DIN1(n5556),
    .DIN1_t(n5556_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX5982),
    .Q_t(WX5982_t)
  );


  nor2s3
  U1591
  (
    .DIN1(n5560),
    .DIN1_t(n5560_t),
    .DIN2(n6731),
    .DIN2_t(n6731_t),
    .Q(WX5980),
    .Q_t(WX5980_t)
  );


  nor2s3
  U1592
  (
    .DIN1(n5564),
    .DIN1_t(n5564_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5978),
    .Q_t(WX5978_t)
  );


  nor2s3
  U1593
  (
    .DIN1(n5568),
    .DIN1_t(n5568_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5976),
    .Q_t(WX5976_t)
  );


  and2s3
  U1594
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5572),
    .DIN2_t(n5572_t),
    .Q(WX5974),
    .Q_t(WX5974_t)
  );


  and2s3
  U1595
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5577),
    .DIN2_t(n5577_t),
    .Q(WX5972),
    .Q_t(WX5972_t)
  );


  and2s3
  U1596
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5582),
    .DIN2_t(n5582_t),
    .Q(WX5970),
    .Q_t(WX5970_t)
  );


  and2s3
  U1597
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5587),
    .DIN2_t(n5587_t),
    .Q(WX5968),
    .Q_t(WX5968_t)
  );


  and2s3
  U1598
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5592),
    .DIN2_t(n5592_t),
    .Q(WX5966),
    .Q_t(WX5966_t)
  );


  and2s3
  U1599
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5597),
    .DIN2_t(n5597_t),
    .Q(WX5964),
    .Q_t(WX5964_t)
  );


  and2s3
  U1600
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5602),
    .DIN2_t(n5602_t),
    .Q(WX5962),
    .Q_t(WX5962_t)
  );


  and2s3
  U1601
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5607),
    .DIN2_t(n5607_t),
    .Q(WX5960),
    .Q_t(WX5960_t)
  );


  and2s3
  U1602
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5612),
    .DIN2_t(n5612_t),
    .Q(WX5958),
    .Q_t(WX5958_t)
  );


  and2s3
  U1603
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5617),
    .DIN2_t(n5617_t),
    .Q(WX5956),
    .Q_t(WX5956_t)
  );


  and2s3
  U1604
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5622),
    .DIN2_t(n5622_t),
    .Q(WX5954),
    .Q_t(WX5954_t)
  );


  and2s3
  U1605
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5627),
    .DIN2_t(n5627_t),
    .Q(WX5952),
    .Q_t(WX5952_t)
  );


  and2s3
  U1606
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5632),
    .DIN2_t(n5632_t),
    .Q(WX5950),
    .Q_t(WX5950_t)
  );


  and2s3
  U1607
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5637),
    .DIN2_t(n5637_t),
    .Q(WX5948),
    .Q_t(WX5948_t)
  );


  and2s3
  U1608
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5642),
    .DIN2_t(n5642_t),
    .Q(WX5946),
    .Q_t(WX5946_t)
  );


  and2s3
  U1609
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5647),
    .DIN2_t(n5647_t),
    .Q(WX5944),
    .Q_t(WX5944_t)
  );


  and2s3
  U1610
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5507),
    .DIN2_t(n5507_t),
    .Q(WX5942),
    .Q_t(WX5942_t)
  );


  and2s3
  U1611
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5511),
    .DIN2_t(n5511_t),
    .Q(WX5940),
    .Q_t(WX5940_t)
  );


  and2s3
  U1612
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5515),
    .DIN2_t(n5515_t),
    .Q(WX5938),
    .Q_t(WX5938_t)
  );


  and2s3
  U1613
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5519),
    .DIN2_t(n5519_t),
    .Q(WX5936),
    .Q_t(WX5936_t)
  );


  and2s3
  U1614
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5523),
    .DIN2_t(n5523_t),
    .Q(WX5934),
    .Q_t(WX5934_t)
  );


  and2s3
  U1615
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5527),
    .DIN2_t(n5527_t),
    .Q(WX5932),
    .Q_t(WX5932_t)
  );


  and2s3
  U1616
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5531),
    .DIN2_t(n5531_t),
    .Q(WX5930),
    .Q_t(WX5930_t)
  );


  and2s3
  U1617
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5535),
    .DIN2_t(n5535_t),
    .Q(WX5928),
    .Q_t(WX5928_t)
  );


  and2s3
  U1618
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5539),
    .DIN2_t(n5539_t),
    .Q(WX5926),
    .Q_t(WX5926_t)
  );


  and2s3
  U1619
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5543),
    .DIN2_t(n5543_t),
    .Q(WX5924),
    .Q_t(WX5924_t)
  );


  and2s3
  U1620
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5547),
    .DIN2_t(n5547_t),
    .Q(WX5922),
    .Q_t(WX5922_t)
  );


  and2s3
  U1621
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5551),
    .DIN2_t(n5551_t),
    .Q(WX5920),
    .Q_t(WX5920_t)
  );


  and2s3
  U1622
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5555),
    .DIN2_t(n5555_t),
    .Q(WX5918),
    .Q_t(WX5918_t)
  );


  and2s3
  U1623
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5559),
    .DIN2_t(n5559_t),
    .Q(WX5916),
    .Q_t(WX5916_t)
  );


  and2s3
  U1624
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5563),
    .DIN2_t(n5563_t),
    .Q(WX5914),
    .Q_t(WX5914_t)
  );


  and2s3
  U1625
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5567),
    .DIN2_t(n5567_t),
    .Q(WX5912),
    .Q_t(WX5912_t)
  );


  nor2s3
  U1626
  (
    .DIN1(n5571),
    .DIN1_t(n5571_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5910),
    .Q_t(WX5910_t)
  );


  nor2s3
  U1627
  (
    .DIN1(n5576),
    .DIN1_t(n5576_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5908),
    .Q_t(WX5908_t)
  );


  nor2s3
  U1628
  (
    .DIN1(n5581),
    .DIN1_t(n5581_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5906),
    .Q_t(WX5906_t)
  );


  nor2s3
  U1629
  (
    .DIN1(n5586),
    .DIN1_t(n5586_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5904),
    .Q_t(WX5904_t)
  );


  nor2s3
  U1630
  (
    .DIN1(n5591),
    .DIN1_t(n5591_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5902),
    .Q_t(WX5902_t)
  );


  nor2s3
  U1631
  (
    .DIN1(n5596),
    .DIN1_t(n5596_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5900),
    .Q_t(WX5900_t)
  );


  nor2s3
  U1632
  (
    .DIN1(n5601),
    .DIN1_t(n5601_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5898),
    .Q_t(WX5898_t)
  );


  nor2s3
  U1633
  (
    .DIN1(n5606),
    .DIN1_t(n5606_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5896),
    .Q_t(WX5896_t)
  );


  nor2s3
  U1634
  (
    .DIN1(n5611),
    .DIN1_t(n5611_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5894),
    .Q_t(WX5894_t)
  );


  nor2s3
  U1635
  (
    .DIN1(n5616),
    .DIN1_t(n5616_t),
    .DIN2(n6730),
    .DIN2_t(n6730_t),
    .Q(WX5892),
    .Q_t(WX5892_t)
  );


  nor2s3
  U1636
  (
    .DIN1(n5621),
    .DIN1_t(n5621_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5890),
    .Q_t(WX5890_t)
  );


  nor2s3
  U1637
  (
    .DIN1(n5626),
    .DIN1_t(n5626_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5888),
    .Q_t(WX5888_t)
  );


  nor2s3
  U1638
  (
    .DIN1(n5631),
    .DIN1_t(n5631_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5886),
    .Q_t(WX5886_t)
  );


  nor2s3
  U1639
  (
    .DIN1(n5636),
    .DIN1_t(n5636_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5884),
    .Q_t(WX5884_t)
  );


  nor2s3
  U1640
  (
    .DIN1(n5641),
    .DIN1_t(n5641_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5882),
    .Q_t(WX5882_t)
  );


  nor2s3
  U1641
  (
    .DIN1(n5646),
    .DIN1_t(n5646_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5880),
    .Q_t(WX5880_t)
  );


  nnd4s2
  U1642
  (
    .DIN1(n3409),
    .DIN1_t(n3409_t),
    .DIN2(n3410),
    .DIN2_t(n3410_t),
    .DIN3(n3411),
    .DIN3_t(n3411_t),
    .DIN4(n3412),
    .DIN4_t(n3412_t),
    .Q(WX5878),
    .Q_t(WX5878_t)
  );


  nnd2s3
  U1643
  (
    .DIN1(n2820),
    .DIN1_t(n2820_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3412),
    .Q_t(n3412_t)
  );


  xor2s3
  U1644
  (
    .DIN1(n3413),
    .DIN1_t(n3413_t),
    .DIN2(n3414),
    .DIN2_t(n3414_t),
    .Q(n2820),
    .Q_t(n2820_t)
  );


  xor2s3
  U1645
  (
    .DIN1(n5331),
    .DIN1_t(n5331_t),
    .DIN2(n5332),
    .DIN2_t(n5332_t),
    .Q(n3414),
    .Q_t(n3414_t)
  );


  xnr2s3
  U1646
  (
    .DIN1(n3237),
    .DIN1_t(n3237_t),
    .DIN2(n5333),
    .DIN2_t(n5333_t),
    .Q(n3413),
    .Q_t(n3413_t)
  );


  nnd2s3
  U1647
  (
    .DIN1(n3415),
    .DIN1_t(n3415_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3411),
    .Q_t(n3411_t)
  );


  nnd2s3
  U1648
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2017),
    .DIN2_t(n2017_t),
    .Q(n3410),
    .Q_t(n3410_t)
  );


  nnd2s3
  U1649
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2016),
    .DIN2_t(n2016_t),
    .Q(n3409),
    .Q_t(n3409_t)
  );


  nnd4s2
  U1650
  (
    .DIN1(n3416),
    .DIN1_t(n3416_t),
    .DIN2(n3417),
    .DIN2_t(n3417_t),
    .DIN3(n3418),
    .DIN3_t(n3418_t),
    .DIN4(n3419),
    .DIN4_t(n3419_t),
    .Q(WX5876),
    .Q_t(WX5876_t)
  );


  nnd2s3
  U1651
  (
    .DIN1(n2827),
    .DIN1_t(n2827_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3419),
    .Q_t(n3419_t)
  );


  xor2s3
  U1652
  (
    .DIN1(n3420),
    .DIN1_t(n3420_t),
    .DIN2(n3421),
    .DIN2_t(n3421_t),
    .Q(n2827),
    .Q_t(n2827_t)
  );


  xor2s3
  U1653
  (
    .DIN1(n5335),
    .DIN1_t(n5335_t),
    .DIN2(n5336),
    .DIN2_t(n5336_t),
    .Q(n3421),
    .Q_t(n3421_t)
  );


  xnr2s3
  U1654
  (
    .DIN1(n3238),
    .DIN1_t(n3238_t),
    .DIN2(n5337),
    .DIN2_t(n5337_t),
    .Q(n3420),
    .Q_t(n3420_t)
  );


  nnd2s3
  U1655
  (
    .DIN1(n3422),
    .DIN1_t(n3422_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3418),
    .Q_t(n3418_t)
  );


  nnd2s3
  U1656
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2018),
    .DIN2_t(n2018_t),
    .Q(n3417),
    .Q_t(n3417_t)
  );


  nnd2s3
  U1657
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2015),
    .DIN2_t(n2015_t),
    .Q(n3416),
    .Q_t(n3416_t)
  );


  nnd4s2
  U1658
  (
    .DIN1(n3423),
    .DIN1_t(n3423_t),
    .DIN2(n3424),
    .DIN2_t(n3424_t),
    .DIN3(n3425),
    .DIN3_t(n3425_t),
    .DIN4(n3426),
    .DIN4_t(n3426_t),
    .Q(WX5874),
    .Q_t(WX5874_t)
  );


  nnd2s3
  U1659
  (
    .DIN1(n2834),
    .DIN1_t(n2834_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3426),
    .Q_t(n3426_t)
  );


  xor2s3
  U1660
  (
    .DIN1(n3427),
    .DIN1_t(n3427_t),
    .DIN2(n3428),
    .DIN2_t(n3428_t),
    .Q(n2834),
    .Q_t(n2834_t)
  );


  xor2s3
  U1661
  (
    .DIN1(n5339),
    .DIN1_t(n5339_t),
    .DIN2(n5340),
    .DIN2_t(n5340_t),
    .Q(n3428),
    .Q_t(n3428_t)
  );


  xnr2s3
  U1662
  (
    .DIN1(n3239),
    .DIN1_t(n3239_t),
    .DIN2(n5341),
    .DIN2_t(n5341_t),
    .Q(n3427),
    .Q_t(n3427_t)
  );


  nnd2s3
  U1663
  (
    .DIN1(n3429),
    .DIN1_t(n3429_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3425),
    .Q_t(n3425_t)
  );


  nnd2s3
  U1664
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2019),
    .DIN2_t(n2019_t),
    .Q(n3424),
    .Q_t(n3424_t)
  );


  nnd2s3
  U1665
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2014),
    .DIN2_t(n2014_t),
    .Q(n3423),
    .Q_t(n3423_t)
  );


  nnd4s2
  U1666
  (
    .DIN1(n3430),
    .DIN1_t(n3430_t),
    .DIN2(n3431),
    .DIN2_t(n3431_t),
    .DIN3(n3432),
    .DIN3_t(n3432_t),
    .DIN4(n3433),
    .DIN4_t(n3433_t),
    .Q(WX5872),
    .Q_t(WX5872_t)
  );


  nnd2s3
  U1667
  (
    .DIN1(n2841),
    .DIN1_t(n2841_t),
    .DIN2(n6626),
    .DIN2_t(n6626_t),
    .Q(n3433),
    .Q_t(n3433_t)
  );


  xor2s3
  U1668
  (
    .DIN1(n3434),
    .DIN1_t(n3434_t),
    .DIN2(n3435),
    .DIN2_t(n3435_t),
    .Q(n2841),
    .Q_t(n2841_t)
  );


  xor2s3
  U1669
  (
    .DIN1(n5343),
    .DIN1_t(n5343_t),
    .DIN2(n5344),
    .DIN2_t(n5344_t),
    .Q(n3435),
    .Q_t(n3435_t)
  );


  xnr2s3
  U1670
  (
    .DIN1(n3240),
    .DIN1_t(n3240_t),
    .DIN2(n5345),
    .DIN2_t(n5345_t),
    .Q(n3434),
    .Q_t(n3434_t)
  );


  nnd2s3
  U1671
  (
    .DIN1(n3436),
    .DIN1_t(n3436_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3432),
    .Q_t(n3432_t)
  );


  nnd2s3
  U1672
  (
    .DIN1(n6606),
    .DIN1_t(n6606_t),
    .DIN2(n2020),
    .DIN2_t(n2020_t),
    .Q(n3431),
    .Q_t(n3431_t)
  );


  nnd2s3
  U1673
  (
    .DIN1(n6575),
    .DIN1_t(n6575_t),
    .DIN2(n2013),
    .DIN2_t(n2013_t),
    .Q(n3430),
    .Q_t(n3430_t)
  );


  nnd4s2
  U1674
  (
    .DIN1(n3437),
    .DIN1_t(n3437_t),
    .DIN2(n3438),
    .DIN2_t(n3438_t),
    .DIN3(n3439),
    .DIN3_t(n3439_t),
    .DIN4(n3440),
    .DIN4_t(n3440_t),
    .Q(WX5870),
    .Q_t(WX5870_t)
  );


  nnd2s3
  U1675
  (
    .DIN1(n2848),
    .DIN1_t(n2848_t),
    .DIN2(n6625),
    .DIN2_t(n6625_t),
    .Q(n3440),
    .Q_t(n3440_t)
  );


  xor2s3
  U1676
  (
    .DIN1(n3441),
    .DIN1_t(n3441_t),
    .DIN2(n3442),
    .DIN2_t(n3442_t),
    .Q(n2848),
    .Q_t(n2848_t)
  );


  xor2s3
  U1677
  (
    .DIN1(n5347),
    .DIN1_t(n5347_t),
    .DIN2(n5348),
    .DIN2_t(n5348_t),
    .Q(n3442),
    .Q_t(n3442_t)
  );


  xnr2s3
  U1678
  (
    .DIN1(n3241),
    .DIN1_t(n3241_t),
    .DIN2(n5349),
    .DIN2_t(n5349_t),
    .Q(n3441),
    .Q_t(n3441_t)
  );


  nnd2s3
  U1679
  (
    .DIN1(n3443),
    .DIN1_t(n3443_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3439),
    .Q_t(n3439_t)
  );


  nnd2s3
  U1680
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2021),
    .DIN2_t(n2021_t),
    .Q(n3438),
    .Q_t(n3438_t)
  );


  nnd2s3
  U1681
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2012),
    .DIN2_t(n2012_t),
    .Q(n3437),
    .Q_t(n3437_t)
  );


  nnd4s2
  U1682
  (
    .DIN1(n3444),
    .DIN1_t(n3444_t),
    .DIN2(n3445),
    .DIN2_t(n3445_t),
    .DIN3(n3446),
    .DIN3_t(n3446_t),
    .DIN4(n3447),
    .DIN4_t(n3447_t),
    .Q(WX5868),
    .Q_t(WX5868_t)
  );


  nnd2s3
  U1683
  (
    .DIN1(n2855),
    .DIN1_t(n2855_t),
    .DIN2(n6625),
    .DIN2_t(n6625_t),
    .Q(n3447),
    .Q_t(n3447_t)
  );


  xor2s3
  U1684
  (
    .DIN1(n3448),
    .DIN1_t(n3448_t),
    .DIN2(n3449),
    .DIN2_t(n3449_t),
    .Q(n2855),
    .Q_t(n2855_t)
  );


  xor2s3
  U1685
  (
    .DIN1(n5351),
    .DIN1_t(n5351_t),
    .DIN2(n5352),
    .DIN2_t(n5352_t),
    .Q(n3449),
    .Q_t(n3449_t)
  );


  xnr2s3
  U1686
  (
    .DIN1(n3242),
    .DIN1_t(n3242_t),
    .DIN2(n5353),
    .DIN2_t(n5353_t),
    .Q(n3448),
    .Q_t(n3448_t)
  );


  nnd2s3
  U1687
  (
    .DIN1(n3450),
    .DIN1_t(n3450_t),
    .DIN2(n6658),
    .DIN2_t(n6658_t),
    .Q(n3446),
    .Q_t(n3446_t)
  );


  nnd2s3
  U1688
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2022),
    .DIN2_t(n2022_t),
    .Q(n3445),
    .Q_t(n3445_t)
  );


  nnd2s3
  U1689
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2011),
    .DIN2_t(n2011_t),
    .Q(n3444),
    .Q_t(n3444_t)
  );


  nnd4s2
  U1690
  (
    .DIN1(n3451),
    .DIN1_t(n3451_t),
    .DIN2(n3452),
    .DIN2_t(n3452_t),
    .DIN3(n3453),
    .DIN3_t(n3453_t),
    .DIN4(n3454),
    .DIN4_t(n3454_t),
    .Q(WX5866),
    .Q_t(WX5866_t)
  );


  nnd2s3
  U1691
  (
    .DIN1(n2862),
    .DIN1_t(n2862_t),
    .DIN2(n6625),
    .DIN2_t(n6625_t),
    .Q(n3454),
    .Q_t(n3454_t)
  );


  xor2s3
  U1692
  (
    .DIN1(n3455),
    .DIN1_t(n3455_t),
    .DIN2(n3456),
    .DIN2_t(n3456_t),
    .Q(n2862),
    .Q_t(n2862_t)
  );


  xor2s3
  U1693
  (
    .DIN1(n5355),
    .DIN1_t(n5355_t),
    .DIN2(n5356),
    .DIN2_t(n5356_t),
    .Q(n3456),
    .Q_t(n3456_t)
  );


  xnr2s3
  U1694
  (
    .DIN1(n3243),
    .DIN1_t(n3243_t),
    .DIN2(n5357),
    .DIN2_t(n5357_t),
    .Q(n3455),
    .Q_t(n3455_t)
  );


  nnd2s3
  U1695
  (
    .DIN1(n3457),
    .DIN1_t(n3457_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3453),
    .Q_t(n3453_t)
  );


  nnd2s3
  U1696
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2023),
    .DIN2_t(n2023_t),
    .Q(n3452),
    .Q_t(n3452_t)
  );


  nnd2s3
  U1697
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2010),
    .DIN2_t(n2010_t),
    .Q(n3451),
    .Q_t(n3451_t)
  );


  nnd4s2
  U1698
  (
    .DIN1(n3458),
    .DIN1_t(n3458_t),
    .DIN2(n3459),
    .DIN2_t(n3459_t),
    .DIN3(n3460),
    .DIN3_t(n3460_t),
    .DIN4(n3461),
    .DIN4_t(n3461_t),
    .Q(WX5864),
    .Q_t(WX5864_t)
  );


  nnd2s3
  U1699
  (
    .DIN1(n2869),
    .DIN1_t(n2869_t),
    .DIN2(n6628),
    .DIN2_t(n6628_t),
    .Q(n3461),
    .Q_t(n3461_t)
  );


  xor2s3
  U1700
  (
    .DIN1(n3462),
    .DIN1_t(n3462_t),
    .DIN2(n3463),
    .DIN2_t(n3463_t),
    .Q(n2869),
    .Q_t(n2869_t)
  );


  xor2s3
  U1701
  (
    .DIN1(n5359),
    .DIN1_t(n5359_t),
    .DIN2(n5360),
    .DIN2_t(n5360_t),
    .Q(n3463),
    .Q_t(n3463_t)
  );


  xnr2s3
  U1702
  (
    .DIN1(n3244),
    .DIN1_t(n3244_t),
    .DIN2(n5361),
    .DIN2_t(n5361_t),
    .Q(n3462),
    .Q_t(n3462_t)
  );


  nnd2s3
  U1703
  (
    .DIN1(n3464),
    .DIN1_t(n3464_t),
    .DIN2(n6658),
    .DIN2_t(n6658_t),
    .Q(n3460),
    .Q_t(n3460_t)
  );


  nnd2s3
  U1704
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2024),
    .DIN2_t(n2024_t),
    .Q(n3459),
    .Q_t(n3459_t)
  );


  nnd2s3
  U1705
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2009),
    .DIN2_t(n2009_t),
    .Q(n3458),
    .Q_t(n3458_t)
  );


  nnd4s2
  U1706
  (
    .DIN1(n3465),
    .DIN1_t(n3465_t),
    .DIN2(n3466),
    .DIN2_t(n3466_t),
    .DIN3(n3467),
    .DIN3_t(n3467_t),
    .DIN4(n3468),
    .DIN4_t(n3468_t),
    .Q(WX5862),
    .Q_t(WX5862_t)
  );


  nnd2s3
  U1707
  (
    .DIN1(n2876),
    .DIN1_t(n2876_t),
    .DIN2(n6625),
    .DIN2_t(n6625_t),
    .Q(n3468),
    .Q_t(n3468_t)
  );


  xor2s3
  U1708
  (
    .DIN1(n3469),
    .DIN1_t(n3469_t),
    .DIN2(n3470),
    .DIN2_t(n3470_t),
    .Q(n2876),
    .Q_t(n2876_t)
  );


  xor2s3
  U1709
  (
    .DIN1(n5363),
    .DIN1_t(n5363_t),
    .DIN2(n5364),
    .DIN2_t(n5364_t),
    .Q(n3470),
    .Q_t(n3470_t)
  );


  xnr2s3
  U1710
  (
    .DIN1(n3245),
    .DIN1_t(n3245_t),
    .DIN2(n5365),
    .DIN2_t(n5365_t),
    .Q(n3469),
    .Q_t(n3469_t)
  );


  nnd2s3
  U1711
  (
    .DIN1(n3471),
    .DIN1_t(n3471_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n3467),
    .Q_t(n3467_t)
  );


  nnd2s3
  U1712
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2025),
    .DIN2_t(n2025_t),
    .Q(n3466),
    .Q_t(n3466_t)
  );


  nnd2s3
  U1713
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2008),
    .DIN2_t(n2008_t),
    .Q(n3465),
    .Q_t(n3465_t)
  );


  nnd4s2
  U1714
  (
    .DIN1(n3472),
    .DIN1_t(n3472_t),
    .DIN2(n3473),
    .DIN2_t(n3473_t),
    .DIN3(n3474),
    .DIN3_t(n3474_t),
    .DIN4(n3475),
    .DIN4_t(n3475_t),
    .Q(WX5860),
    .Q_t(WX5860_t)
  );


  nnd2s3
  U1715
  (
    .DIN1(n2883),
    .DIN1_t(n2883_t),
    .DIN2(n6625),
    .DIN2_t(n6625_t),
    .Q(n3475),
    .Q_t(n3475_t)
  );


  xor2s3
  U1716
  (
    .DIN1(n3476),
    .DIN1_t(n3476_t),
    .DIN2(n3477),
    .DIN2_t(n3477_t),
    .Q(n2883),
    .Q_t(n2883_t)
  );


  xor2s3
  U1717
  (
    .DIN1(n5367),
    .DIN1_t(n5367_t),
    .DIN2(n5368),
    .DIN2_t(n5368_t),
    .Q(n3477),
    .Q_t(n3477_t)
  );


  xnr2s3
  U1718
  (
    .DIN1(n3246),
    .DIN1_t(n3246_t),
    .DIN2(n5369),
    .DIN2_t(n5369_t),
    .Q(n3476),
    .Q_t(n3476_t)
  );


  nnd2s3
  U1719
  (
    .DIN1(n3478),
    .DIN1_t(n3478_t),
    .DIN2(n6658),
    .DIN2_t(n6658_t),
    .Q(n3474),
    .Q_t(n3474_t)
  );


  nnd2s3
  U1720
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2026),
    .DIN2_t(n2026_t),
    .Q(n3473),
    .Q_t(n3473_t)
  );


  nnd2s3
  U1721
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2007),
    .DIN2_t(n2007_t),
    .Q(n3472),
    .Q_t(n3472_t)
  );


  nnd4s2
  U1722
  (
    .DIN1(n3479),
    .DIN1_t(n3479_t),
    .DIN2(n3480),
    .DIN2_t(n3480_t),
    .DIN3(n3481),
    .DIN3_t(n3481_t),
    .DIN4(n3482),
    .DIN4_t(n3482_t),
    .Q(WX5858),
    .Q_t(WX5858_t)
  );


  nnd2s3
  U1723
  (
    .DIN1(n2890),
    .DIN1_t(n2890_t),
    .DIN2(n6625),
    .DIN2_t(n6625_t),
    .Q(n3482),
    .Q_t(n3482_t)
  );


  xor2s3
  U1724
  (
    .DIN1(n3483),
    .DIN1_t(n3483_t),
    .DIN2(n3484),
    .DIN2_t(n3484_t),
    .Q(n2890),
    .Q_t(n2890_t)
  );


  xor2s3
  U1725
  (
    .DIN1(n5371),
    .DIN1_t(n5371_t),
    .DIN2(n5372),
    .DIN2_t(n5372_t),
    .Q(n3484),
    .Q_t(n3484_t)
  );


  xnr2s3
  U1726
  (
    .DIN1(n3247),
    .DIN1_t(n3247_t),
    .DIN2(n5373),
    .DIN2_t(n5373_t),
    .Q(n3483),
    .Q_t(n3483_t)
  );


  nnd2s3
  U1727
  (
    .DIN1(n3485),
    .DIN1_t(n3485_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3481),
    .Q_t(n3481_t)
  );


  nnd2s3
  U1728
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2027),
    .DIN2_t(n2027_t),
    .Q(n3480),
    .Q_t(n3480_t)
  );


  nnd2s3
  U1729
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2006),
    .DIN2_t(n2006_t),
    .Q(n3479),
    .Q_t(n3479_t)
  );


  nnd4s2
  U1730
  (
    .DIN1(n3486),
    .DIN1_t(n3486_t),
    .DIN2(n3487),
    .DIN2_t(n3487_t),
    .DIN3(n3488),
    .DIN3_t(n3488_t),
    .DIN4(n3489),
    .DIN4_t(n3489_t),
    .Q(WX5856),
    .Q_t(WX5856_t)
  );


  nnd2s3
  U1731
  (
    .DIN1(n2897),
    .DIN1_t(n2897_t),
    .DIN2(n6625),
    .DIN2_t(n6625_t),
    .Q(n3489),
    .Q_t(n3489_t)
  );


  xor2s3
  U1732
  (
    .DIN1(n3490),
    .DIN1_t(n3490_t),
    .DIN2(n3491),
    .DIN2_t(n3491_t),
    .Q(n2897),
    .Q_t(n2897_t)
  );


  xor2s3
  U1733
  (
    .DIN1(n5375),
    .DIN1_t(n5375_t),
    .DIN2(n5376),
    .DIN2_t(n5376_t),
    .Q(n3491),
    .Q_t(n3491_t)
  );


  xnr2s3
  U1734
  (
    .DIN1(n3248),
    .DIN1_t(n3248_t),
    .DIN2(n5377),
    .DIN2_t(n5377_t),
    .Q(n3490),
    .Q_t(n3490_t)
  );


  nnd2s3
  U1735
  (
    .DIN1(n3492),
    .DIN1_t(n3492_t),
    .DIN2(n6658),
    .DIN2_t(n6658_t),
    .Q(n3488),
    .Q_t(n3488_t)
  );


  nnd2s3
  U1736
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2028),
    .DIN2_t(n2028_t),
    .Q(n3487),
    .Q_t(n3487_t)
  );


  nnd2s3
  U1737
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2005),
    .DIN2_t(n2005_t),
    .Q(n3486),
    .Q_t(n3486_t)
  );


  nnd4s2
  U1738
  (
    .DIN1(n3493),
    .DIN1_t(n3493_t),
    .DIN2(n3494),
    .DIN2_t(n3494_t),
    .DIN3(n3495),
    .DIN3_t(n3495_t),
    .DIN4(n3496),
    .DIN4_t(n3496_t),
    .Q(WX5854),
    .Q_t(WX5854_t)
  );


  nnd2s3
  U1739
  (
    .DIN1(n2904),
    .DIN1_t(n2904_t),
    .DIN2(n6625),
    .DIN2_t(n6625_t),
    .Q(n3496),
    .Q_t(n3496_t)
  );


  xor2s3
  U1740
  (
    .DIN1(n3497),
    .DIN1_t(n3497_t),
    .DIN2(n3498),
    .DIN2_t(n3498_t),
    .Q(n2904),
    .Q_t(n2904_t)
  );


  xor2s3
  U1741
  (
    .DIN1(n5379),
    .DIN1_t(n5379_t),
    .DIN2(n5380),
    .DIN2_t(n5380_t),
    .Q(n3498),
    .Q_t(n3498_t)
  );


  xnr2s3
  U1742
  (
    .DIN1(n3249),
    .DIN1_t(n3249_t),
    .DIN2(n5381),
    .DIN2_t(n5381_t),
    .Q(n3497),
    .Q_t(n3497_t)
  );


  nnd2s3
  U1743
  (
    .DIN1(n3499),
    .DIN1_t(n3499_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3495),
    .Q_t(n3495_t)
  );


  nnd2s3
  U1744
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2029),
    .DIN2_t(n2029_t),
    .Q(n3494),
    .Q_t(n3494_t)
  );


  nnd2s3
  U1745
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2004),
    .DIN2_t(n2004_t),
    .Q(n3493),
    .Q_t(n3493_t)
  );


  nnd4s2
  U1746
  (
    .DIN1(n3500),
    .DIN1_t(n3500_t),
    .DIN2(n3501),
    .DIN2_t(n3501_t),
    .DIN3(n3502),
    .DIN3_t(n3502_t),
    .DIN4(n3503),
    .DIN4_t(n3503_t),
    .Q(WX5852),
    .Q_t(WX5852_t)
  );


  nnd2s3
  U1747
  (
    .DIN1(n2911),
    .DIN1_t(n2911_t),
    .DIN2(n6625),
    .DIN2_t(n6625_t),
    .Q(n3503),
    .Q_t(n3503_t)
  );


  xor2s3
  U1748
  (
    .DIN1(n3504),
    .DIN1_t(n3504_t),
    .DIN2(n3505),
    .DIN2_t(n3505_t),
    .Q(n2911),
    .Q_t(n2911_t)
  );


  xor2s3
  U1749
  (
    .DIN1(n5383),
    .DIN1_t(n5383_t),
    .DIN2(n5384),
    .DIN2_t(n5384_t),
    .Q(n3505),
    .Q_t(n3505_t)
  );


  xnr2s3
  U1750
  (
    .DIN1(n3250),
    .DIN1_t(n3250_t),
    .DIN2(n5385),
    .DIN2_t(n5385_t),
    .Q(n3504),
    .Q_t(n3504_t)
  );


  nnd2s3
  U1751
  (
    .DIN1(n3506),
    .DIN1_t(n3506_t),
    .DIN2(n6658),
    .DIN2_t(n6658_t),
    .Q(n3502),
    .Q_t(n3502_t)
  );


  nnd2s3
  U1752
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2030),
    .DIN2_t(n2030_t),
    .Q(n3501),
    .Q_t(n3501_t)
  );


  nnd2s3
  U1753
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2003),
    .DIN2_t(n2003_t),
    .Q(n3500),
    .Q_t(n3500_t)
  );


  nnd4s2
  U1754
  (
    .DIN1(n3507),
    .DIN1_t(n3507_t),
    .DIN2(n3508),
    .DIN2_t(n3508_t),
    .DIN3(n3509),
    .DIN3_t(n3509_t),
    .DIN4(n3510),
    .DIN4_t(n3510_t),
    .Q(WX5850),
    .Q_t(WX5850_t)
  );


  nnd2s3
  U1755
  (
    .DIN1(n2918),
    .DIN1_t(n2918_t),
    .DIN2(n6625),
    .DIN2_t(n6625_t),
    .Q(n3510),
    .Q_t(n3510_t)
  );


  xor2s3
  U1756
  (
    .DIN1(n3511),
    .DIN1_t(n3511_t),
    .DIN2(n3512),
    .DIN2_t(n3512_t),
    .Q(n2918),
    .Q_t(n2918_t)
  );


  xor2s3
  U1757
  (
    .DIN1(n5387),
    .DIN1_t(n5387_t),
    .DIN2(n5388),
    .DIN2_t(n5388_t),
    .Q(n3512),
    .Q_t(n3512_t)
  );


  xnr2s3
  U1758
  (
    .DIN1(n3251),
    .DIN1_t(n3251_t),
    .DIN2(n5389),
    .DIN2_t(n5389_t),
    .Q(n3511),
    .Q_t(n3511_t)
  );


  nnd2s3
  U1759
  (
    .DIN1(n3513),
    .DIN1_t(n3513_t),
    .DIN2(n6659),
    .DIN2_t(n6659_t),
    .Q(n3509),
    .Q_t(n3509_t)
  );


  nnd2s3
  U1760
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2031),
    .DIN2_t(n2031_t),
    .Q(n3508),
    .Q_t(n3508_t)
  );


  nnd2s3
  U1761
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2002),
    .DIN2_t(n2002_t),
    .Q(n3507),
    .Q_t(n3507_t)
  );


  nnd4s2
  U1762
  (
    .DIN1(n3514),
    .DIN1_t(n3514_t),
    .DIN2(n3515),
    .DIN2_t(n3515_t),
    .DIN3(n3516),
    .DIN3_t(n3516_t),
    .DIN4(n3517),
    .DIN4_t(n3517_t),
    .Q(WX5848),
    .Q_t(WX5848_t)
  );


  nnd2s3
  U1763
  (
    .DIN1(n2925),
    .DIN1_t(n2925_t),
    .DIN2(n6630),
    .DIN2_t(n6630_t),
    .Q(n3517),
    .Q_t(n3517_t)
  );


  xor2s3
  U1764
  (
    .DIN1(n3518),
    .DIN1_t(n3518_t),
    .DIN2(n3519),
    .DIN2_t(n3519_t),
    .Q(n2925),
    .Q_t(n2925_t)
  );


  xor2s3
  U1765
  (
    .DIN1(n5391),
    .DIN1_t(n5391_t),
    .DIN2(n5392),
    .DIN2_t(n5392_t),
    .Q(n3519),
    .Q_t(n3519_t)
  );


  xnr2s3
  U1766
  (
    .DIN1(n3252),
    .DIN1_t(n3252_t),
    .DIN2(n5393),
    .DIN2_t(n5393_t),
    .Q(n3518),
    .Q_t(n3518_t)
  );


  nnd2s3
  U1767
  (
    .DIN1(n3520),
    .DIN1_t(n3520_t),
    .DIN2(n6658),
    .DIN2_t(n6658_t),
    .Q(n3516),
    .Q_t(n3516_t)
  );


  nnd2s3
  U1768
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2032),
    .DIN2_t(n2032_t),
    .Q(n3515),
    .Q_t(n3515_t)
  );


  nnd2s3
  U1769
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2001),
    .DIN2_t(n2001_t),
    .Q(n3514),
    .Q_t(n3514_t)
  );


  nnd4s2
  U1770
  (
    .DIN1(n3521),
    .DIN1_t(n3521_t),
    .DIN2(n3522),
    .DIN2_t(n3522_t),
    .DIN3(n3523),
    .DIN3_t(n3523_t),
    .DIN4(n3524),
    .DIN4_t(n3524_t),
    .Q(WX5846),
    .Q_t(WX5846_t)
  );


  nnd2s3
  U1771
  (
    .DIN1(n2933),
    .DIN1_t(n2933_t),
    .DIN2(n6647),
    .DIN2_t(n6647_t),
    .Q(n3524),
    .Q_t(n3524_t)
  );


  xor2s3
  U1772
  (
    .DIN1(n3525),
    .DIN1_t(n3525_t),
    .DIN2(n3526),
    .DIN2_t(n3526_t),
    .Q(n2933),
    .Q_t(n2933_t)
  );


  xor2s3
  U1773
  (
    .DIN1(n5397),
    .DIN1_t(n5397_t),
    .DIN2(n3527),
    .DIN2_t(n3527_t),
    .Q(n3526),
    .Q_t(n3526_t)
  );


  xor2s3
  U1774
  (
    .DIN1(n5395),
    .DIN1_t(n5395_t),
    .DIN2(n5396),
    .DIN2_t(n5396_t),
    .Q(n3527),
    .Q_t(n3527_t)
  );


  xor2s3
  U1775
  (
    .DIN1(n5398),
    .DIN1_t(n5398_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3525),
    .Q_t(n3525_t)
  );


  nnd2s3
  U1776
  (
    .DIN1(n3528),
    .DIN1_t(n3528_t),
    .DIN2(n6678),
    .DIN2_t(n6678_t),
    .Q(n3523),
    .Q_t(n3523_t)
  );


  nnd2s3
  U1777
  (
    .DIN1(n6605),
    .DIN1_t(n6605_t),
    .DIN2(n2033),
    .DIN2_t(n2033_t),
    .Q(n3522),
    .Q_t(n3522_t)
  );


  nnd2s3
  U1778
  (
    .DIN1(n6574),
    .DIN1_t(n6574_t),
    .DIN2(n2000),
    .DIN2_t(n2000_t),
    .Q(n3521),
    .Q_t(n3521_t)
  );


  nnd4s2
  U1779
  (
    .DIN1(n3529),
    .DIN1_t(n3529_t),
    .DIN2(n3530),
    .DIN2_t(n3530_t),
    .DIN3(n3531),
    .DIN3_t(n3531_t),
    .DIN4(n3532),
    .DIN4_t(n3532_t),
    .Q(WX5844),
    .Q_t(WX5844_t)
  );


  nnd2s3
  U1780
  (
    .DIN1(n2941),
    .DIN1_t(n2941_t),
    .DIN2(n6647),
    .DIN2_t(n6647_t),
    .Q(n3532),
    .Q_t(n3532_t)
  );


  xor2s3
  U1781
  (
    .DIN1(n3533),
    .DIN1_t(n3533_t),
    .DIN2(n3534),
    .DIN2_t(n3534_t),
    .Q(n2941),
    .Q_t(n2941_t)
  );


  xor2s3
  U1782
  (
    .DIN1(n5402),
    .DIN1_t(n5402_t),
    .DIN2(n3535),
    .DIN2_t(n3535_t),
    .Q(n3534),
    .Q_t(n3534_t)
  );


  xor2s3
  U1783
  (
    .DIN1(n5400),
    .DIN1_t(n5400_t),
    .DIN2(n5401),
    .DIN2_t(n5401_t),
    .Q(n3535),
    .Q_t(n3535_t)
  );


  xor2s3
  U1784
  (
    .DIN1(n5403),
    .DIN1_t(n5403_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3533),
    .Q_t(n3533_t)
  );


  nnd2s3
  U1785
  (
    .DIN1(n3536),
    .DIN1_t(n3536_t),
    .DIN2(n6678),
    .DIN2_t(n6678_t),
    .Q(n3531),
    .Q_t(n3531_t)
  );


  nnd2s3
  U1786
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2034),
    .DIN2_t(n2034_t),
    .Q(n3530),
    .Q_t(n3530_t)
  );


  nnd2s3
  U1787
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1999),
    .DIN2_t(n1999_t),
    .Q(n3529),
    .Q_t(n3529_t)
  );


  nnd4s2
  U1788
  (
    .DIN1(n3537),
    .DIN1_t(n3537_t),
    .DIN2(n3538),
    .DIN2_t(n3538_t),
    .DIN3(n3539),
    .DIN3_t(n3539_t),
    .DIN4(n3540),
    .DIN4_t(n3540_t),
    .Q(WX5842),
    .Q_t(WX5842_t)
  );


  nnd2s3
  U1789
  (
    .DIN1(n2949),
    .DIN1_t(n2949_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3540),
    .Q_t(n3540_t)
  );


  xor2s3
  U1790
  (
    .DIN1(n3541),
    .DIN1_t(n3541_t),
    .DIN2(n3542),
    .DIN2_t(n3542_t),
    .Q(n2949),
    .Q_t(n2949_t)
  );


  xor2s3
  U1791
  (
    .DIN1(n5407),
    .DIN1_t(n5407_t),
    .DIN2(n3543),
    .DIN2_t(n3543_t),
    .Q(n3542),
    .Q_t(n3542_t)
  );


  xor2s3
  U1792
  (
    .DIN1(n5405),
    .DIN1_t(n5405_t),
    .DIN2(n5406),
    .DIN2_t(n5406_t),
    .Q(n3543),
    .Q_t(n3543_t)
  );


  xor2s3
  U1793
  (
    .DIN1(n5408),
    .DIN1_t(n5408_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3541),
    .Q_t(n3541_t)
  );


  nnd2s3
  U1794
  (
    .DIN1(n3544),
    .DIN1_t(n3544_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3539),
    .Q_t(n3539_t)
  );


  nnd2s3
  U1795
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2035),
    .DIN2_t(n2035_t),
    .Q(n3538),
    .Q_t(n3538_t)
  );


  nnd2s3
  U1796
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1998),
    .DIN2_t(n1998_t),
    .Q(n3537),
    .Q_t(n3537_t)
  );


  nnd4s2
  U1797
  (
    .DIN1(n3545),
    .DIN1_t(n3545_t),
    .DIN2(n3546),
    .DIN2_t(n3546_t),
    .DIN3(n3547),
    .DIN3_t(n3547_t),
    .DIN4(n3548),
    .DIN4_t(n3548_t),
    .Q(WX5840),
    .Q_t(WX5840_t)
  );


  nnd2s3
  U1798
  (
    .DIN1(n2957),
    .DIN1_t(n2957_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3548),
    .Q_t(n3548_t)
  );


  xor2s3
  U1799
  (
    .DIN1(n3549),
    .DIN1_t(n3549_t),
    .DIN2(n3550),
    .DIN2_t(n3550_t),
    .Q(n2957),
    .Q_t(n2957_t)
  );


  xor2s3
  U1800
  (
    .DIN1(n5412),
    .DIN1_t(n5412_t),
    .DIN2(n3551),
    .DIN2_t(n3551_t),
    .Q(n3550),
    .Q_t(n3550_t)
  );


  xor2s3
  U1801
  (
    .DIN1(n5410),
    .DIN1_t(n5410_t),
    .DIN2(n5411),
    .DIN2_t(n5411_t),
    .Q(n3551),
    .Q_t(n3551_t)
  );


  xor2s3
  U1802
  (
    .DIN1(n5413),
    .DIN1_t(n5413_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3549),
    .Q_t(n3549_t)
  );


  nnd2s3
  U1803
  (
    .DIN1(n3552),
    .DIN1_t(n3552_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3547),
    .Q_t(n3547_t)
  );


  nnd2s3
  U1804
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2036),
    .DIN2_t(n2036_t),
    .Q(n3546),
    .Q_t(n3546_t)
  );


  nnd2s3
  U1805
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1997),
    .DIN2_t(n1997_t),
    .Q(n3545),
    .Q_t(n3545_t)
  );


  nnd4s2
  U1806
  (
    .DIN1(n3553),
    .DIN1_t(n3553_t),
    .DIN2(n3554),
    .DIN2_t(n3554_t),
    .DIN3(n3555),
    .DIN3_t(n3555_t),
    .DIN4(n3556),
    .DIN4_t(n3556_t),
    .Q(WX5838),
    .Q_t(WX5838_t)
  );


  nnd2s3
  U1807
  (
    .DIN1(n2965),
    .DIN1_t(n2965_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3556),
    .Q_t(n3556_t)
  );


  xor2s3
  U1808
  (
    .DIN1(n3557),
    .DIN1_t(n3557_t),
    .DIN2(n3558),
    .DIN2_t(n3558_t),
    .Q(n2965),
    .Q_t(n2965_t)
  );


  xor2s3
  U1809
  (
    .DIN1(n5417),
    .DIN1_t(n5417_t),
    .DIN2(n3559),
    .DIN2_t(n3559_t),
    .Q(n3558),
    .Q_t(n3558_t)
  );


  xor2s3
  U1810
  (
    .DIN1(n5415),
    .DIN1_t(n5415_t),
    .DIN2(n5416),
    .DIN2_t(n5416_t),
    .Q(n3559),
    .Q_t(n3559_t)
  );


  xor2s3
  U1811
  (
    .DIN1(n5418),
    .DIN1_t(n5418_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3557),
    .Q_t(n3557_t)
  );


  nnd2s3
  U1812
  (
    .DIN1(n3560),
    .DIN1_t(n3560_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3555),
    .Q_t(n3555_t)
  );


  nnd2s3
  U1813
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2037),
    .DIN2_t(n2037_t),
    .Q(n3554),
    .Q_t(n3554_t)
  );


  nnd2s3
  U1814
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1996),
    .DIN2_t(n1996_t),
    .Q(n3553),
    .Q_t(n3553_t)
  );


  nnd4s2
  U1815
  (
    .DIN1(n3561),
    .DIN1_t(n3561_t),
    .DIN2(n3562),
    .DIN2_t(n3562_t),
    .DIN3(n3563),
    .DIN3_t(n3563_t),
    .DIN4(n3564),
    .DIN4_t(n3564_t),
    .Q(WX5836),
    .Q_t(WX5836_t)
  );


  nnd2s3
  U1816
  (
    .DIN1(n2973),
    .DIN1_t(n2973_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3564),
    .Q_t(n3564_t)
  );


  xor2s3
  U1817
  (
    .DIN1(n3565),
    .DIN1_t(n3565_t),
    .DIN2(n3566),
    .DIN2_t(n3566_t),
    .Q(n2973),
    .Q_t(n2973_t)
  );


  xor2s3
  U1818
  (
    .DIN1(n5422),
    .DIN1_t(n5422_t),
    .DIN2(n3567),
    .DIN2_t(n3567_t),
    .Q(n3566),
    .Q_t(n3566_t)
  );


  xor2s3
  U1819
  (
    .DIN1(n5420),
    .DIN1_t(n5420_t),
    .DIN2(n5421),
    .DIN2_t(n5421_t),
    .Q(n3567),
    .Q_t(n3567_t)
  );


  xor2s3
  U1820
  (
    .DIN1(n5423),
    .DIN1_t(n5423_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3565),
    .Q_t(n3565_t)
  );


  nnd2s3
  U1821
  (
    .DIN1(n3568),
    .DIN1_t(n3568_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3563),
    .Q_t(n3563_t)
  );


  nnd2s3
  U1822
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2038),
    .DIN2_t(n2038_t),
    .Q(n3562),
    .Q_t(n3562_t)
  );


  nnd2s3
  U1823
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1995),
    .DIN2_t(n1995_t),
    .Q(n3561),
    .Q_t(n3561_t)
  );


  nnd4s2
  U1824
  (
    .DIN1(n3569),
    .DIN1_t(n3569_t),
    .DIN2(n3570),
    .DIN2_t(n3570_t),
    .DIN3(n3571),
    .DIN3_t(n3571_t),
    .DIN4(n3572),
    .DIN4_t(n3572_t),
    .Q(WX5834),
    .Q_t(WX5834_t)
  );


  nnd2s3
  U1825
  (
    .DIN1(n2981),
    .DIN1_t(n2981_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3572),
    .Q_t(n3572_t)
  );


  xor2s3
  U1826
  (
    .DIN1(n3573),
    .DIN1_t(n3573_t),
    .DIN2(n3574),
    .DIN2_t(n3574_t),
    .Q(n2981),
    .Q_t(n2981_t)
  );


  xor2s3
  U1827
  (
    .DIN1(n5427),
    .DIN1_t(n5427_t),
    .DIN2(n3575),
    .DIN2_t(n3575_t),
    .Q(n3574),
    .Q_t(n3574_t)
  );


  xor2s3
  U1828
  (
    .DIN1(n5425),
    .DIN1_t(n5425_t),
    .DIN2(n5426),
    .DIN2_t(n5426_t),
    .Q(n3575),
    .Q_t(n3575_t)
  );


  xor2s3
  U1829
  (
    .DIN1(n5428),
    .DIN1_t(n5428_t),
    .DIN2(n6689),
    .DIN2_t(n6689_t),
    .Q(n3573),
    .Q_t(n3573_t)
  );


  nnd2s3
  U1830
  (
    .DIN1(n3576),
    .DIN1_t(n3576_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3571),
    .Q_t(n3571_t)
  );


  nnd2s3
  U1831
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2039),
    .DIN2_t(n2039_t),
    .Q(n3570),
    .Q_t(n3570_t)
  );


  nnd2s3
  U1832
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1994),
    .DIN2_t(n1994_t),
    .Q(n3569),
    .Q_t(n3569_t)
  );


  nnd4s2
  U1833
  (
    .DIN1(n3577),
    .DIN1_t(n3577_t),
    .DIN2(n3578),
    .DIN2_t(n3578_t),
    .DIN3(n3579),
    .DIN3_t(n3579_t),
    .DIN4(n3580),
    .DIN4_t(n3580_t),
    .Q(WX5832),
    .Q_t(WX5832_t)
  );


  nnd2s3
  U1834
  (
    .DIN1(n2989),
    .DIN1_t(n2989_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3580),
    .Q_t(n3580_t)
  );


  xor2s3
  U1835
  (
    .DIN1(n3581),
    .DIN1_t(n3581_t),
    .DIN2(n3582),
    .DIN2_t(n3582_t),
    .Q(n2989),
    .Q_t(n2989_t)
  );


  xor2s3
  U1836
  (
    .DIN1(n5432),
    .DIN1_t(n5432_t),
    .DIN2(n3583),
    .DIN2_t(n3583_t),
    .Q(n3582),
    .Q_t(n3582_t)
  );


  xor2s3
  U1837
  (
    .DIN1(n5430),
    .DIN1_t(n5430_t),
    .DIN2(n5431),
    .DIN2_t(n5431_t),
    .Q(n3583),
    .Q_t(n3583_t)
  );


  xor2s3
  U1838
  (
    .DIN1(n5433),
    .DIN1_t(n5433_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3581),
    .Q_t(n3581_t)
  );


  nnd2s3
  U1839
  (
    .DIN1(n3584),
    .DIN1_t(n3584_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3579),
    .Q_t(n3579_t)
  );


  nnd2s3
  U1840
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2040),
    .DIN2_t(n2040_t),
    .Q(n3578),
    .Q_t(n3578_t)
  );


  nnd2s3
  U1841
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1993),
    .DIN2_t(n1993_t),
    .Q(n3577),
    .Q_t(n3577_t)
  );


  nnd4s2
  U1842
  (
    .DIN1(n3585),
    .DIN1_t(n3585_t),
    .DIN2(n3586),
    .DIN2_t(n3586_t),
    .DIN3(n3587),
    .DIN3_t(n3587_t),
    .DIN4(n3588),
    .DIN4_t(n3588_t),
    .Q(WX5830),
    .Q_t(WX5830_t)
  );


  nnd2s3
  U1843
  (
    .DIN1(n2997),
    .DIN1_t(n2997_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3588),
    .Q_t(n3588_t)
  );


  xor2s3
  U1844
  (
    .DIN1(n3589),
    .DIN1_t(n3589_t),
    .DIN2(n3590),
    .DIN2_t(n3590_t),
    .Q(n2997),
    .Q_t(n2997_t)
  );


  xor2s3
  U1845
  (
    .DIN1(n5437),
    .DIN1_t(n5437_t),
    .DIN2(n3591),
    .DIN2_t(n3591_t),
    .Q(n3590),
    .Q_t(n3590_t)
  );


  xor2s3
  U1846
  (
    .DIN1(n5435),
    .DIN1_t(n5435_t),
    .DIN2(n5436),
    .DIN2_t(n5436_t),
    .Q(n3591),
    .Q_t(n3591_t)
  );


  xor2s3
  U1847
  (
    .DIN1(n5438),
    .DIN1_t(n5438_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3589),
    .Q_t(n3589_t)
  );


  nnd2s3
  U1848
  (
    .DIN1(n3592),
    .DIN1_t(n3592_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3587),
    .Q_t(n3587_t)
  );


  nnd2s3
  U1849
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2041),
    .DIN2_t(n2041_t),
    .Q(n3586),
    .Q_t(n3586_t)
  );


  nnd2s3
  U1850
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1992),
    .DIN2_t(n1992_t),
    .Q(n3585),
    .Q_t(n3585_t)
  );


  nnd4s2
  U1851
  (
    .DIN1(n3593),
    .DIN1_t(n3593_t),
    .DIN2(n3594),
    .DIN2_t(n3594_t),
    .DIN3(n3595),
    .DIN3_t(n3595_t),
    .DIN4(n3596),
    .DIN4_t(n3596_t),
    .Q(WX5828),
    .Q_t(WX5828_t)
  );


  nnd2s3
  U1852
  (
    .DIN1(n3005),
    .DIN1_t(n3005_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3596),
    .Q_t(n3596_t)
  );


  xor2s3
  U1853
  (
    .DIN1(n3597),
    .DIN1_t(n3597_t),
    .DIN2(n3598),
    .DIN2_t(n3598_t),
    .Q(n3005),
    .Q_t(n3005_t)
  );


  xor2s3
  U1854
  (
    .DIN1(n5442),
    .DIN1_t(n5442_t),
    .DIN2(n3599),
    .DIN2_t(n3599_t),
    .Q(n3598),
    .Q_t(n3598_t)
  );


  xor2s3
  U1855
  (
    .DIN1(n5440),
    .DIN1_t(n5440_t),
    .DIN2(n5441),
    .DIN2_t(n5441_t),
    .Q(n3599),
    .Q_t(n3599_t)
  );


  xor2s3
  U1856
  (
    .DIN1(n5443),
    .DIN1_t(n5443_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3597),
    .Q_t(n3597_t)
  );


  nnd2s3
  U1857
  (
    .DIN1(n3600),
    .DIN1_t(n3600_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3595),
    .Q_t(n3595_t)
  );


  nnd2s3
  U1858
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2042),
    .DIN2_t(n2042_t),
    .Q(n3594),
    .Q_t(n3594_t)
  );


  nnd2s3
  U1859
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1991),
    .DIN2_t(n1991_t),
    .Q(n3593),
    .Q_t(n3593_t)
  );


  nnd4s2
  U1860
  (
    .DIN1(n3601),
    .DIN1_t(n3601_t),
    .DIN2(n3602),
    .DIN2_t(n3602_t),
    .DIN3(n3603),
    .DIN3_t(n3603_t),
    .DIN4(n3604),
    .DIN4_t(n3604_t),
    .Q(WX5826),
    .Q_t(WX5826_t)
  );


  nnd2s3
  U1861
  (
    .DIN1(n3013),
    .DIN1_t(n3013_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3604),
    .Q_t(n3604_t)
  );


  xor2s3
  U1862
  (
    .DIN1(n3605),
    .DIN1_t(n3605_t),
    .DIN2(n3606),
    .DIN2_t(n3606_t),
    .Q(n3013),
    .Q_t(n3013_t)
  );


  xor2s3
  U1863
  (
    .DIN1(n5447),
    .DIN1_t(n5447_t),
    .DIN2(n3607),
    .DIN2_t(n3607_t),
    .Q(n3606),
    .Q_t(n3606_t)
  );


  xor2s3
  U1864
  (
    .DIN1(n5445),
    .DIN1_t(n5445_t),
    .DIN2(n5446),
    .DIN2_t(n5446_t),
    .Q(n3607),
    .Q_t(n3607_t)
  );


  xor2s3
  U1865
  (
    .DIN1(n5448),
    .DIN1_t(n5448_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3605),
    .Q_t(n3605_t)
  );


  nnd2s3
  U1866
  (
    .DIN1(n3608),
    .DIN1_t(n3608_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3603),
    .Q_t(n3603_t)
  );


  nnd2s3
  U1867
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2043),
    .DIN2_t(n2043_t),
    .Q(n3602),
    .Q_t(n3602_t)
  );


  nnd2s3
  U1868
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1990),
    .DIN2_t(n1990_t),
    .Q(n3601),
    .Q_t(n3601_t)
  );


  nnd4s2
  U1869
  (
    .DIN1(n3609),
    .DIN1_t(n3609_t),
    .DIN2(n3610),
    .DIN2_t(n3610_t),
    .DIN3(n3611),
    .DIN3_t(n3611_t),
    .DIN4(n3612),
    .DIN4_t(n3612_t),
    .Q(WX5824),
    .Q_t(WX5824_t)
  );


  nnd2s3
  U1870
  (
    .DIN1(n3021),
    .DIN1_t(n3021_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3612),
    .Q_t(n3612_t)
  );


  xor2s3
  U1871
  (
    .DIN1(n3613),
    .DIN1_t(n3613_t),
    .DIN2(n3614),
    .DIN2_t(n3614_t),
    .Q(n3021),
    .Q_t(n3021_t)
  );


  xor2s3
  U1872
  (
    .DIN1(n5452),
    .DIN1_t(n5452_t),
    .DIN2(n3615),
    .DIN2_t(n3615_t),
    .Q(n3614),
    .Q_t(n3614_t)
  );


  xor2s3
  U1873
  (
    .DIN1(n5450),
    .DIN1_t(n5450_t),
    .DIN2(n5451),
    .DIN2_t(n5451_t),
    .Q(n3615),
    .Q_t(n3615_t)
  );


  xor2s3
  U1874
  (
    .DIN1(n5453),
    .DIN1_t(n5453_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3613),
    .Q_t(n3613_t)
  );


  nnd2s3
  U1875
  (
    .DIN1(n3616),
    .DIN1_t(n3616_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3611),
    .Q_t(n3611_t)
  );


  nnd2s3
  U1876
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2044),
    .DIN2_t(n2044_t),
    .Q(n3610),
    .Q_t(n3610_t)
  );


  nnd2s3
  U1877
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1989),
    .DIN2_t(n1989_t),
    .Q(n3609),
    .Q_t(n3609_t)
  );


  nnd4s2
  U1878
  (
    .DIN1(n3617),
    .DIN1_t(n3617_t),
    .DIN2(n3618),
    .DIN2_t(n3618_t),
    .DIN3(n3619),
    .DIN3_t(n3619_t),
    .DIN4(n3620),
    .DIN4_t(n3620_t),
    .Q(WX5822),
    .Q_t(WX5822_t)
  );


  nnd2s3
  U1879
  (
    .DIN1(n3029),
    .DIN1_t(n3029_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3620),
    .Q_t(n3620_t)
  );


  xor2s3
  U1880
  (
    .DIN1(n3621),
    .DIN1_t(n3621_t),
    .DIN2(n3622),
    .DIN2_t(n3622_t),
    .Q(n3029),
    .Q_t(n3029_t)
  );


  xor2s3
  U1881
  (
    .DIN1(n5457),
    .DIN1_t(n5457_t),
    .DIN2(n3623),
    .DIN2_t(n3623_t),
    .Q(n3622),
    .Q_t(n3622_t)
  );


  xor2s3
  U1882
  (
    .DIN1(n5455),
    .DIN1_t(n5455_t),
    .DIN2(n5456),
    .DIN2_t(n5456_t),
    .Q(n3623),
    .Q_t(n3623_t)
  );


  xor2s3
  U1883
  (
    .DIN1(n5458),
    .DIN1_t(n5458_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3621),
    .Q_t(n3621_t)
  );


  nnd2s3
  U1884
  (
    .DIN1(n3624),
    .DIN1_t(n3624_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3619),
    .Q_t(n3619_t)
  );


  nnd2s3
  U1885
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2045),
    .DIN2_t(n2045_t),
    .Q(n3618),
    .Q_t(n3618_t)
  );


  nnd2s3
  U1886
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1988),
    .DIN2_t(n1988_t),
    .Q(n3617),
    .Q_t(n3617_t)
  );


  nnd4s2
  U1887
  (
    .DIN1(n3625),
    .DIN1_t(n3625_t),
    .DIN2(n3626),
    .DIN2_t(n3626_t),
    .DIN3(n3627),
    .DIN3_t(n3627_t),
    .DIN4(n3628),
    .DIN4_t(n3628_t),
    .Q(WX5820),
    .Q_t(WX5820_t)
  );


  nnd2s3
  U1888
  (
    .DIN1(n3037),
    .DIN1_t(n3037_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3628),
    .Q_t(n3628_t)
  );


  xor2s3
  U1889
  (
    .DIN1(n3629),
    .DIN1_t(n3629_t),
    .DIN2(n3630),
    .DIN2_t(n3630_t),
    .Q(n3037),
    .Q_t(n3037_t)
  );


  xor2s3
  U1890
  (
    .DIN1(n5462),
    .DIN1_t(n5462_t),
    .DIN2(n3631),
    .DIN2_t(n3631_t),
    .Q(n3630),
    .Q_t(n3630_t)
  );


  xor2s3
  U1891
  (
    .DIN1(n5460),
    .DIN1_t(n5460_t),
    .DIN2(n5461),
    .DIN2_t(n5461_t),
    .Q(n3631),
    .Q_t(n3631_t)
  );


  xor2s3
  U1892
  (
    .DIN1(n5463),
    .DIN1_t(n5463_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3629),
    .Q_t(n3629_t)
  );


  nnd2s3
  U1893
  (
    .DIN1(n3632),
    .DIN1_t(n3632_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3627),
    .Q_t(n3627_t)
  );


  nnd2s3
  U1894
  (
    .DIN1(n6604),
    .DIN1_t(n6604_t),
    .DIN2(n2046),
    .DIN2_t(n2046_t),
    .Q(n3626),
    .Q_t(n3626_t)
  );


  nnd2s3
  U1895
  (
    .DIN1(n6573),
    .DIN1_t(n6573_t),
    .DIN2(n1987),
    .DIN2_t(n1987_t),
    .Q(n3625),
    .Q_t(n3625_t)
  );


  nnd4s2
  U1896
  (
    .DIN1(n3633),
    .DIN1_t(n3633_t),
    .DIN2(n3634),
    .DIN2_t(n3634_t),
    .DIN3(n3635),
    .DIN3_t(n3635_t),
    .DIN4(n3636),
    .DIN4_t(n3636_t),
    .Q(WX5818),
    .Q_t(WX5818_t)
  );


  nnd2s3
  U1897
  (
    .DIN1(n3045),
    .DIN1_t(n3045_t),
    .DIN2(n6646),
    .DIN2_t(n6646_t),
    .Q(n3636),
    .Q_t(n3636_t)
  );


  xor2s3
  U1898
  (
    .DIN1(n3637),
    .DIN1_t(n3637_t),
    .DIN2(n3638),
    .DIN2_t(n3638_t),
    .Q(n3045),
    .Q_t(n3045_t)
  );


  xor2s3
  U1899
  (
    .DIN1(n5467),
    .DIN1_t(n5467_t),
    .DIN2(n3639),
    .DIN2_t(n3639_t),
    .Q(n3638),
    .Q_t(n3638_t)
  );


  xor2s3
  U1900
  (
    .DIN1(n5465),
    .DIN1_t(n5465_t),
    .DIN2(n5466),
    .DIN2_t(n5466_t),
    .Q(n3639),
    .Q_t(n3639_t)
  );


  xor2s3
  U1901
  (
    .DIN1(n5468),
    .DIN1_t(n5468_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3637),
    .Q_t(n3637_t)
  );


  nnd2s3
  U1902
  (
    .DIN1(n3640),
    .DIN1_t(n3640_t),
    .DIN2(n6677),
    .DIN2_t(n6677_t),
    .Q(n3635),
    .Q_t(n3635_t)
  );


  nnd2s3
  U1903
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2047),
    .DIN2_t(n2047_t),
    .Q(n3634),
    .Q_t(n3634_t)
  );


  nnd2s3
  U1904
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n1986),
    .DIN2_t(n1986_t),
    .Q(n3633),
    .Q_t(n3633_t)
  );


  nnd4s2
  U1905
  (
    .DIN1(n3641),
    .DIN1_t(n3641_t),
    .DIN2(n3642),
    .DIN2_t(n3642_t),
    .DIN3(n3643),
    .DIN3_t(n3643_t),
    .DIN4(n3644),
    .DIN4_t(n3644_t),
    .Q(WX5816),
    .Q_t(WX5816_t)
  );


  nnd2s3
  U1906
  (
    .DIN1(n3053),
    .DIN1_t(n3053_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3644),
    .Q_t(n3644_t)
  );


  xor2s3
  U1907
  (
    .DIN1(n3645),
    .DIN1_t(n3645_t),
    .DIN2(n3646),
    .DIN2_t(n3646_t),
    .Q(n3053),
    .Q_t(n3053_t)
  );


  xor2s3
  U1908
  (
    .DIN1(n5472),
    .DIN1_t(n5472_t),
    .DIN2(n3647),
    .DIN2_t(n3647_t),
    .Q(n3646),
    .Q_t(n3646_t)
  );


  xor2s3
  U1909
  (
    .DIN1(n5470),
    .DIN1_t(n5470_t),
    .DIN2(n5471),
    .DIN2_t(n5471_t),
    .Q(n3647),
    .Q_t(n3647_t)
  );


  xor2s3
  U1910
  (
    .DIN1(n5473),
    .DIN1_t(n5473_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3645),
    .Q_t(n3645_t)
  );


  nnd2s3
  U1911
  (
    .DIN1(n3648),
    .DIN1_t(n3648_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3643),
    .Q_t(n3643_t)
  );


  nnd2s3
  U1912
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2048),
    .DIN2_t(n2048_t),
    .Q(n3642),
    .Q_t(n3642_t)
  );


  nnd2s3
  U1913
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n1985),
    .DIN2_t(n1985_t),
    .Q(n3641),
    .Q_t(n3641_t)
  );


  nor2s3
  U1914
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n2048),
    .DIN2_t(n2048_t),
    .Q(WX5718),
    .Q_t(WX5718_t)
  );


  nor2s3
  U1915
  (
    .DIN1(n5476),
    .DIN1_t(n5476_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5716),
    .Q_t(WX5716_t)
  );


  nor2s3
  U1916
  (
    .DIN1(n5477),
    .DIN1_t(n5477_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5714),
    .Q_t(WX5714_t)
  );


  nor2s3
  U1917
  (
    .DIN1(n5478),
    .DIN1_t(n5478_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5712),
    .Q_t(WX5712_t)
  );


  nor2s3
  U1918
  (
    .DIN1(n5479),
    .DIN1_t(n5479_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5710),
    .Q_t(WX5710_t)
  );


  nor2s3
  U1919
  (
    .DIN1(n5480),
    .DIN1_t(n5480_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5708),
    .Q_t(WX5708_t)
  );


  nor2s3
  U1920
  (
    .DIN1(n5481),
    .DIN1_t(n5481_t),
    .DIN2(n6729),
    .DIN2_t(n6729_t),
    .Q(WX5706),
    .Q_t(WX5706_t)
  );


  nor2s3
  U1921
  (
    .DIN1(n5482),
    .DIN1_t(n5482_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX5704),
    .Q_t(WX5704_t)
  );


  nor2s3
  U1922
  (
    .DIN1(n5483),
    .DIN1_t(n5483_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX5702),
    .Q_t(WX5702_t)
  );


  nor2s3
  U1923
  (
    .DIN1(n5484),
    .DIN1_t(n5484_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX5700),
    .Q_t(WX5700_t)
  );


  nor2s3
  U1924
  (
    .DIN1(n5485),
    .DIN1_t(n5485_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX5698),
    .Q_t(WX5698_t)
  );


  nor2s3
  U1925
  (
    .DIN1(n5486),
    .DIN1_t(n5486_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX5696),
    .Q_t(WX5696_t)
  );


  nor2s3
  U1926
  (
    .DIN1(n5487),
    .DIN1_t(n5487_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX5694),
    .Q_t(WX5694_t)
  );


  nor2s3
  U1927
  (
    .DIN1(n5488),
    .DIN1_t(n5488_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX5692),
    .Q_t(WX5692_t)
  );


  nor2s3
  U1928
  (
    .DIN1(n5489),
    .DIN1_t(n5489_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX5690),
    .Q_t(WX5690_t)
  );


  nor2s3
  U1929
  (
    .DIN1(n5490),
    .DIN1_t(n5490_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX5688),
    .Q_t(WX5688_t)
  );


  nor2s3
  U1930
  (
    .DIN1(n5491),
    .DIN1_t(n5491_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX5686),
    .Q_t(WX5686_t)
  );


  nor2s3
  U1931
  (
    .DIN1(n5492),
    .DIN1_t(n5492_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX5684),
    .Q_t(WX5684_t)
  );


  nor2s3
  U1932
  (
    .DIN1(n5493),
    .DIN1_t(n5493_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5682),
    .Q_t(WX5682_t)
  );


  nor2s3
  U1933
  (
    .DIN1(n5494),
    .DIN1_t(n5494_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5680),
    .Q_t(WX5680_t)
  );


  nor2s3
  U1934
  (
    .DIN1(n5495),
    .DIN1_t(n5495_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5678),
    .Q_t(WX5678_t)
  );


  nor2s3
  U1935
  (
    .DIN1(n5496),
    .DIN1_t(n5496_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5676),
    .Q_t(WX5676_t)
  );


  nor2s3
  U1936
  (
    .DIN1(n5497),
    .DIN1_t(n5497_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5674),
    .Q_t(WX5674_t)
  );


  nor2s3
  U1937
  (
    .DIN1(n5498),
    .DIN1_t(n5498_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5672),
    .Q_t(WX5672_t)
  );


  nor2s3
  U1938
  (
    .DIN1(n5499),
    .DIN1_t(n5499_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5670),
    .Q_t(WX5670_t)
  );


  nor2s3
  U1939
  (
    .DIN1(n5500),
    .DIN1_t(n5500_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5668),
    .Q_t(WX5668_t)
  );


  nor2s3
  U1940
  (
    .DIN1(n5501),
    .DIN1_t(n5501_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5666),
    .Q_t(WX5666_t)
  );


  nor2s3
  U1941
  (
    .DIN1(n5502),
    .DIN1_t(n5502_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5664),
    .Q_t(WX5664_t)
  );


  nor2s3
  U1942
  (
    .DIN1(n5503),
    .DIN1_t(n5503_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5662),
    .Q_t(WX5662_t)
  );


  nor2s3
  U1943
  (
    .DIN1(n5504),
    .DIN1_t(n5504_t),
    .DIN2(n6727),
    .DIN2_t(n6727_t),
    .Q(WX5660),
    .Q_t(WX5660_t)
  );


  nor2s3
  U1944
  (
    .DIN1(n5505),
    .DIN1_t(n5505_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX5658),
    .Q_t(WX5658_t)
  );


  nor2s3
  U1945
  (
    .DIN1(n5506),
    .DIN1_t(n5506_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX5656),
    .Q_t(WX5656_t)
  );


  nor2s3
  U1946
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n2304),
    .DIN2_t(n2304_t),
    .Q(WX546),
    .Q_t(WX546_t)
  );


  nor2s3
  U1947
  (
    .DIN1(n6179),
    .DIN1_t(n6179_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX544),
    .Q_t(WX544_t)
  );


  nor2s3
  U1948
  (
    .DIN1(n6180),
    .DIN1_t(n6180_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX542),
    .Q_t(WX542_t)
  );


  nor2s3
  U1949
  (
    .DIN1(n6181),
    .DIN1_t(n6181_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX540),
    .Q_t(WX540_t)
  );


  nor2s3
  U1950
  (
    .DIN1(n6182),
    .DIN1_t(n6182_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX538),
    .Q_t(WX538_t)
  );


  nor2s3
  U1951
  (
    .DIN1(n6183),
    .DIN1_t(n6183_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX536),
    .Q_t(WX536_t)
  );


  nor2s3
  U1952
  (
    .DIN1(n6184),
    .DIN1_t(n6184_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX534),
    .Q_t(WX534_t)
  );


  nor2s3
  U1953
  (
    .DIN1(n6185),
    .DIN1_t(n6185_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX532),
    .Q_t(WX532_t)
  );


  nor2s3
  U1954
  (
    .DIN1(n6186),
    .DIN1_t(n6186_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX530),
    .Q_t(WX530_t)
  );


  nor2s3
  U1955
  (
    .DIN1(n6187),
    .DIN1_t(n6187_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX528),
    .Q_t(WX528_t)
  );


  nor2s3
  U1956
  (
    .DIN1(n6188),
    .DIN1_t(n6188_t),
    .DIN2(n6726),
    .DIN2_t(n6726_t),
    .Q(WX526),
    .Q_t(WX526_t)
  );


  nor2s3
  U1957
  (
    .DIN1(n6189),
    .DIN1_t(n6189_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX524),
    .Q_t(WX524_t)
  );


  nor2s3
  U1958
  (
    .DIN1(n6190),
    .DIN1_t(n6190_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX522),
    .Q_t(WX522_t)
  );


  nor2s3
  U1959
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n3649),
    .DIN2_t(n3649_t),
    .Q(WX5205),
    .Q_t(WX5205_t)
  );


  xor2s3
  U1960
  (
    .DIN1(n5645),
    .DIN1_t(n5645_t),
    .DIN2(n5825),
    .DIN2_t(n5825_t),
    .Q(n3649),
    .Q_t(n3649_t)
  );


  nor2s3
  U1961
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n3650),
    .DIN2_t(n3650_t),
    .Q(WX5203),
    .Q_t(WX5203_t)
  );


  xor2s3
  U1962
  (
    .DIN1(n5640),
    .DIN1_t(n5640_t),
    .DIN2(n5820),
    .DIN2_t(n5820_t),
    .Q(n3650),
    .Q_t(n3650_t)
  );


  nor2s3
  U1963
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n3651),
    .DIN2_t(n3651_t),
    .Q(WX5201),
    .Q_t(WX5201_t)
  );


  xor2s3
  U1964
  (
    .DIN1(n5635),
    .DIN1_t(n5635_t),
    .DIN2(n5815),
    .DIN2_t(n5815_t),
    .Q(n3651),
    .Q_t(n3651_t)
  );


  nor2s3
  U1965
  (
    .DIN1(n6191),
    .DIN1_t(n6191_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX520),
    .Q_t(WX520_t)
  );


  nor2s3
  U1966
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n3652),
    .DIN2_t(n3652_t),
    .Q(WX5199),
    .Q_t(WX5199_t)
  );


  xor2s3
  U1967
  (
    .DIN1(n5630),
    .DIN1_t(n5630_t),
    .DIN2(n5810),
    .DIN2_t(n5810_t),
    .Q(n3652),
    .Q_t(n3652_t)
  );


  nor2s3
  U1968
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n3653),
    .DIN2_t(n3653_t),
    .Q(WX5197),
    .Q_t(WX5197_t)
  );


  xor2s3
  U1969
  (
    .DIN1(n5625),
    .DIN1_t(n5625_t),
    .DIN2(n5805),
    .DIN2_t(n5805_t),
    .Q(n3653),
    .Q_t(n3653_t)
  );


  nor2s3
  U1970
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n3654),
    .DIN2_t(n3654_t),
    .Q(WX5195),
    .Q_t(WX5195_t)
  );


  xor2s3
  U1971
  (
    .DIN1(n5620),
    .DIN1_t(n5620_t),
    .DIN2(n5800),
    .DIN2_t(n5800_t),
    .Q(n3654),
    .Q_t(n3654_t)
  );


  nor2s3
  U1972
  (
    .DIN1(n6788),
    .DIN1_t(n6788_t),
    .DIN2(n3655),
    .DIN2_t(n3655_t),
    .Q(WX5193),
    .Q_t(WX5193_t)
  );


  xor2s3
  U1973
  (
    .DIN1(n5615),
    .DIN1_t(n5615_t),
    .DIN2(n5795),
    .DIN2_t(n5795_t),
    .Q(n3655),
    .Q_t(n3655_t)
  );


  nor2s3
  U1974
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n3656),
    .DIN2_t(n3656_t),
    .Q(WX5191),
    .Q_t(WX5191_t)
  );


  xor2s3
  U1975
  (
    .DIN1(n5610),
    .DIN1_t(n5610_t),
    .DIN2(n5790),
    .DIN2_t(n5790_t),
    .Q(n3656),
    .Q_t(n3656_t)
  );


  nor2s3
  U1976
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n3657),
    .DIN2_t(n3657_t),
    .Q(WX5189),
    .Q_t(WX5189_t)
  );


  xor2s3
  U1977
  (
    .DIN1(n5605),
    .DIN1_t(n5605_t),
    .DIN2(n5785),
    .DIN2_t(n5785_t),
    .Q(n3657),
    .Q_t(n3657_t)
  );


  nor2s3
  U1978
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n3658),
    .DIN2_t(n3658_t),
    .Q(WX5187),
    .Q_t(WX5187_t)
  );


  xor2s3
  U1979
  (
    .DIN1(n5600),
    .DIN1_t(n5600_t),
    .DIN2(n5780),
    .DIN2_t(n5780_t),
    .Q(n3658),
    .Q_t(n3658_t)
  );


  nor2s3
  U1980
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n3659),
    .DIN2_t(n3659_t),
    .Q(WX5185),
    .Q_t(WX5185_t)
  );


  xor2s3
  U1981
  (
    .DIN1(n5595),
    .DIN1_t(n5595_t),
    .DIN2(n5775),
    .DIN2_t(n5775_t),
    .Q(n3659),
    .Q_t(n3659_t)
  );


  nor2s3
  U1982
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n3660),
    .DIN2_t(n3660_t),
    .Q(WX5183),
    .Q_t(WX5183_t)
  );


  xor2s3
  U1983
  (
    .DIN1(n5590),
    .DIN1_t(n5590_t),
    .DIN2(n5770),
    .DIN2_t(n5770_t),
    .Q(n3660),
    .Q_t(n3660_t)
  );


  nor2s3
  U1984
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n3661),
    .DIN2_t(n3661_t),
    .Q(WX5181),
    .Q_t(WX5181_t)
  );


  xor2s3
  U1985
  (
    .DIN1(n5585),
    .DIN1_t(n5585_t),
    .DIN2(n5765),
    .DIN2_t(n5765_t),
    .Q(n3661),
    .Q_t(n3661_t)
  );


  nor2s3
  U1986
  (
    .DIN1(n6192),
    .DIN1_t(n6192_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX518),
    .Q_t(WX518_t)
  );


  nor2s3
  U1987
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n3662),
    .DIN2_t(n3662_t),
    .Q(WX5179),
    .Q_t(WX5179_t)
  );


  xor2s3
  U1988
  (
    .DIN1(n5580),
    .DIN1_t(n5580_t),
    .DIN2(n5760),
    .DIN2_t(n5760_t),
    .Q(n3662),
    .Q_t(n3662_t)
  );


  nor2s3
  U1989
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n3663),
    .DIN2_t(n3663_t),
    .Q(WX5177),
    .Q_t(WX5177_t)
  );


  xor2s3
  U1990
  (
    .DIN1(n5575),
    .DIN1_t(n5575_t),
    .DIN2(n5755),
    .DIN2_t(n5755_t),
    .Q(n3663),
    .Q_t(n3663_t)
  );


  nor2s3
  U1991
  (
    .DIN1(n3664),
    .DIN1_t(n3664_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX5175),
    .Q_t(WX5175_t)
  );


  xnr2s3
  U1992
  (
    .DIN1(n5750),
    .DIN1_t(n5750_t),
    .DIN2(n3665),
    .DIN2_t(n3665_t),
    .Q(n3664),
    .Q_t(n3664_t)
  );


  xor2s3
  U1993
  (
    .DIN1(n5570),
    .DIN1_t(n5570_t),
    .DIN2(n5650),
    .DIN2_t(n5650_t),
    .Q(n3665),
    .Q_t(n3665_t)
  );


  nor2s3
  U1994
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n3666),
    .DIN2_t(n3666_t),
    .Q(WX5173),
    .Q_t(WX5173_t)
  );


  xor2s3
  U1995
  (
    .DIN1(n5566),
    .DIN1_t(n5566_t),
    .DIN2(n3284),
    .DIN2_t(n3284_t),
    .Q(n3666),
    .Q_t(n3666_t)
  );


  nor2s3
  U1996
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n3667),
    .DIN2_t(n3667_t),
    .Q(WX5171),
    .Q_t(WX5171_t)
  );


  xor2s3
  U1997
  (
    .DIN1(n5562),
    .DIN1_t(n5562_t),
    .DIN2(n3283),
    .DIN2_t(n3283_t),
    .Q(n3667),
    .Q_t(n3667_t)
  );


  nor2s3
  U1998
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n3668),
    .DIN2_t(n3668_t),
    .Q(WX5169),
    .Q_t(WX5169_t)
  );


  xor2s3
  U1999
  (
    .DIN1(n5558),
    .DIN1_t(n5558_t),
    .DIN2(n3282),
    .DIN2_t(n3282_t),
    .Q(n3668),
    .Q_t(n3668_t)
  );


  nor2s3
  U2000
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n3669),
    .DIN2_t(n3669_t),
    .Q(WX5167),
    .Q_t(WX5167_t)
  );


  xor2s3
  U2001
  (
    .DIN1(n5554),
    .DIN1_t(n5554_t),
    .DIN2(n3281),
    .DIN2_t(n3281_t),
    .Q(n3669),
    .Q_t(n3669_t)
  );


  nor2s3
  U2002
  (
    .DIN1(n3670),
    .DIN1_t(n3670_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX5165),
    .Q_t(WX5165_t)
  );


  xnr2s3
  U2003
  (
    .DIN1(n3280),
    .DIN1_t(n3280_t),
    .DIN2(n3671),
    .DIN2_t(n3671_t),
    .Q(n3670),
    .Q_t(n3670_t)
  );


  xor2s3
  U2004
  (
    .DIN1(n5550),
    .DIN1_t(n5550_t),
    .DIN2(n5650),
    .DIN2_t(n5650_t),
    .Q(n3671),
    .Q_t(n3671_t)
  );


  nor2s3
  U2005
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n3672),
    .DIN2_t(n3672_t),
    .Q(WX5163),
    .Q_t(WX5163_t)
  );


  xor2s3
  U2006
  (
    .DIN1(n5546),
    .DIN1_t(n5546_t),
    .DIN2(n3279),
    .DIN2_t(n3279_t),
    .Q(n3672),
    .Q_t(n3672_t)
  );


  nor2s3
  U2007
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n3673),
    .DIN2_t(n3673_t),
    .Q(WX5161),
    .Q_t(WX5161_t)
  );


  xor2s3
  U2008
  (
    .DIN1(n5542),
    .DIN1_t(n5542_t),
    .DIN2(n3278),
    .DIN2_t(n3278_t),
    .Q(n3673),
    .Q_t(n3673_t)
  );


  nor2s3
  U2009
  (
    .DIN1(n6193),
    .DIN1_t(n6193_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX516),
    .Q_t(WX516_t)
  );


  nor2s3
  U2010
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n3674),
    .DIN2_t(n3674_t),
    .Q(WX5159),
    .Q_t(WX5159_t)
  );


  xor2s3
  U2011
  (
    .DIN1(n5538),
    .DIN1_t(n5538_t),
    .DIN2(n3277),
    .DIN2_t(n3277_t),
    .Q(n3674),
    .Q_t(n3674_t)
  );


  nor2s3
  U2012
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n3675),
    .DIN2_t(n3675_t),
    .Q(WX5157),
    .Q_t(WX5157_t)
  );


  xor2s3
  U2013
  (
    .DIN1(n5534),
    .DIN1_t(n5534_t),
    .DIN2(n3276),
    .DIN2_t(n3276_t),
    .Q(n3675),
    .Q_t(n3675_t)
  );


  nor2s3
  U2014
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n3676),
    .DIN2_t(n3676_t),
    .Q(WX5155),
    .Q_t(WX5155_t)
  );


  xor2s3
  U2015
  (
    .DIN1(n5530),
    .DIN1_t(n5530_t),
    .DIN2(n3275),
    .DIN2_t(n3275_t),
    .Q(n3676),
    .Q_t(n3676_t)
  );


  nor2s3
  U2016
  (
    .DIN1(n6788),
    .DIN1_t(n6788_t),
    .DIN2(n3677),
    .DIN2_t(n3677_t),
    .Q(WX5153),
    .Q_t(WX5153_t)
  );


  xor2s3
  U2017
  (
    .DIN1(n5526),
    .DIN1_t(n5526_t),
    .DIN2(n3274),
    .DIN2_t(n3274_t),
    .Q(n3677),
    .Q_t(n3677_t)
  );


  nor2s3
  U2018
  (
    .DIN1(n3678),
    .DIN1_t(n3678_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX5151),
    .Q_t(WX5151_t)
  );


  xnr2s3
  U2019
  (
    .DIN1(n3273),
    .DIN1_t(n3273_t),
    .DIN2(n3679),
    .DIN2_t(n3679_t),
    .Q(n3678),
    .Q_t(n3678_t)
  );


  xor2s3
  U2020
  (
    .DIN1(n5522),
    .DIN1_t(n5522_t),
    .DIN2(n5650),
    .DIN2_t(n5650_t),
    .Q(n3679),
    .Q_t(n3679_t)
  );


  nor2s3
  U2021
  (
    .DIN1(n6788),
    .DIN1_t(n6788_t),
    .DIN2(n3680),
    .DIN2_t(n3680_t),
    .Q(WX5149),
    .Q_t(WX5149_t)
  );


  xor2s3
  U2022
  (
    .DIN1(n5518),
    .DIN1_t(n5518_t),
    .DIN2(n3272),
    .DIN2_t(n3272_t),
    .Q(n3680),
    .Q_t(n3680_t)
  );


  nor2s3
  U2023
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n3681),
    .DIN2_t(n3681_t),
    .Q(WX5147),
    .Q_t(WX5147_t)
  );


  xor2s3
  U2024
  (
    .DIN1(n5514),
    .DIN1_t(n5514_t),
    .DIN2(n3271),
    .DIN2_t(n3271_t),
    .Q(n3681),
    .Q_t(n3681_t)
  );


  nor2s3
  U2025
  (
    .DIN1(n6788),
    .DIN1_t(n6788_t),
    .DIN2(n3682),
    .DIN2_t(n3682_t),
    .Q(WX5145),
    .Q_t(WX5145_t)
  );


  xor2s3
  U2026
  (
    .DIN1(n5510),
    .DIN1_t(n5510_t),
    .DIN2(n3270),
    .DIN2_t(n3270_t),
    .Q(n3682),
    .Q_t(n3682_t)
  );


  nor2s3
  U2027
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n3683),
    .DIN2_t(n3683_t),
    .Q(WX5143),
    .Q_t(WX5143_t)
  );


  xor2s3
  U2028
  (
    .DIN1(n5650),
    .DIN1_t(n5650_t),
    .DIN2(n3269),
    .DIN2_t(n3269_t),
    .Q(n3683),
    .Q_t(n3683_t)
  );


  nor2s3
  U2029
  (
    .DIN1(n6194),
    .DIN1_t(n6194_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX514),
    .Q_t(WX514_t)
  );


  nor2s3
  U2030
  (
    .DIN1(n6195),
    .DIN1_t(n6195_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX512),
    .Q_t(WX512_t)
  );


  nor2s3
  U2031
  (
    .DIN1(n6196),
    .DIN1_t(n6196_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX510),
    .Q_t(WX510_t)
  );


  nor2s3
  U2032
  (
    .DIN1(n6286),
    .DIN1_t(n6286_t),
    .DIN2(n6725),
    .DIN2_t(n6725_t),
    .Q(WX508),
    .Q_t(WX508_t)
  );


  nor2s3
  U2033
  (
    .DIN1(n6342),
    .DIN1_t(n6342_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX506),
    .Q_t(WX506_t)
  );


  nor2s3
  U2034
  (
    .DIN1(n6354),
    .DIN1_t(n6354_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX504),
    .Q_t(WX504_t)
  );


  nor2s3
  U2035
  (
    .DIN1(n6376),
    .DIN1_t(n6376_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX502),
    .Q_t(WX502_t)
  );


  nor2s3
  U2036
  (
    .DIN1(n6377),
    .DIN1_t(n6377_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX500),
    .Q_t(WX500_t)
  );


  nor2s3
  U2037
  (
    .DIN1(n6378),
    .DIN1_t(n6378_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX498),
    .Q_t(WX498_t)
  );


  nor2s3
  U2038
  (
    .DIN1(n6379),
    .DIN1_t(n6379_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX496),
    .Q_t(WX496_t)
  );


  nor2s3
  U2039
  (
    .DIN1(n6380),
    .DIN1_t(n6380_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX494),
    .Q_t(WX494_t)
  );


  nor2s3
  U2040
  (
    .DIN1(n6381),
    .DIN1_t(n6381_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX492),
    .Q_t(WX492_t)
  );


  nor2s3
  U2041
  (
    .DIN1(n6382),
    .DIN1_t(n6382_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX490),
    .Q_t(WX490_t)
  );


  nor2s3
  U2042
  (
    .DIN1(n6431),
    .DIN1_t(n6431_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX488),
    .Q_t(WX488_t)
  );


  nor2s3
  U2043
  (
    .DIN1(n6432),
    .DIN1_t(n6432_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX486),
    .Q_t(WX486_t)
  );


  nor2s3
  U2044
  (
    .DIN1(n6433),
    .DIN1_t(n6433_t),
    .DIN2(n6724),
    .DIN2_t(n6724_t),
    .Q(WX484),
    .Q_t(WX484_t)
  );


  nor2s3
  U2045
  (
    .DIN1(n5685),
    .DIN1_t(n5685_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX4777),
    .Q_t(WX4777_t)
  );


  nor2s3
  U2046
  (
    .DIN1(n5689),
    .DIN1_t(n5689_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX4775),
    .Q_t(WX4775_t)
  );


  nor2s3
  U2047
  (
    .DIN1(n5693),
    .DIN1_t(n5693_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX4773),
    .Q_t(WX4773_t)
  );


  nor2s3
  U2048
  (
    .DIN1(n5697),
    .DIN1_t(n5697_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX4771),
    .Q_t(WX4771_t)
  );


  nor2s3
  U2049
  (
    .DIN1(n5701),
    .DIN1_t(n5701_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX4769),
    .Q_t(WX4769_t)
  );


  nor2s3
  U2050
  (
    .DIN1(n5705),
    .DIN1_t(n5705_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX4767),
    .Q_t(WX4767_t)
  );


  nor2s3
  U2051
  (
    .DIN1(n5709),
    .DIN1_t(n5709_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX4765),
    .Q_t(WX4765_t)
  );


  nor2s3
  U2052
  (
    .DIN1(n5713),
    .DIN1_t(n5713_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX4763),
    .Q_t(WX4763_t)
  );


  nor2s3
  U2053
  (
    .DIN1(n5717),
    .DIN1_t(n5717_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX4761),
    .Q_t(WX4761_t)
  );


  nor2s3
  U2054
  (
    .DIN1(n5721),
    .DIN1_t(n5721_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX4759),
    .Q_t(WX4759_t)
  );


  nor2s3
  U2055
  (
    .DIN1(n5725),
    .DIN1_t(n5725_t),
    .DIN2(n6723),
    .DIN2_t(n6723_t),
    .Q(WX4757),
    .Q_t(WX4757_t)
  );


  nor2s3
  U2056
  (
    .DIN1(n5729),
    .DIN1_t(n5729_t),
    .DIN2(n6728),
    .DIN2_t(n6728_t),
    .Q(WX4755),
    .Q_t(WX4755_t)
  );


  nor2s3
  U2057
  (
    .DIN1(n5733),
    .DIN1_t(n5733_t),
    .DIN2(n6734),
    .DIN2_t(n6734_t),
    .Q(WX4753),
    .Q_t(WX4753_t)
  );


  nor2s3
  U2058
  (
    .DIN1(n5737),
    .DIN1_t(n5737_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX4751),
    .Q_t(WX4751_t)
  );


  nor2s3
  U2059
  (
    .DIN1(n5741),
    .DIN1_t(n5741_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX4749),
    .Q_t(WX4749_t)
  );


  nor2s3
  U2060
  (
    .DIN1(n5745),
    .DIN1_t(n5745_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX4747),
    .Q_t(WX4747_t)
  );


  nor2s3
  U2061
  (
    .DIN1(n5749),
    .DIN1_t(n5749_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX4745),
    .Q_t(WX4745_t)
  );


  nor2s3
  U2062
  (
    .DIN1(n5754),
    .DIN1_t(n5754_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX4743),
    .Q_t(WX4743_t)
  );


  nor2s3
  U2063
  (
    .DIN1(n5759),
    .DIN1_t(n5759_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX4741),
    .Q_t(WX4741_t)
  );


  nor2s3
  U2064
  (
    .DIN1(n5764),
    .DIN1_t(n5764_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX4739),
    .Q_t(WX4739_t)
  );


  nor2s3
  U2065
  (
    .DIN1(n5769),
    .DIN1_t(n5769_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX4737),
    .Q_t(WX4737_t)
  );


  nor2s3
  U2066
  (
    .DIN1(n5774),
    .DIN1_t(n5774_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX4735),
    .Q_t(WX4735_t)
  );


  nor2s3
  U2067
  (
    .DIN1(n5779),
    .DIN1_t(n5779_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX4733),
    .Q_t(WX4733_t)
  );


  nor2s3
  U2068
  (
    .DIN1(n5784),
    .DIN1_t(n5784_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX4731),
    .Q_t(WX4731_t)
  );


  nor2s3
  U2069
  (
    .DIN1(n5789),
    .DIN1_t(n5789_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX4729),
    .Q_t(WX4729_t)
  );


  nor2s3
  U2070
  (
    .DIN1(n5794),
    .DIN1_t(n5794_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX4727),
    .Q_t(WX4727_t)
  );


  nor2s3
  U2071
  (
    .DIN1(n5799),
    .DIN1_t(n5799_t),
    .DIN2(n6788),
    .DIN2_t(n6788_t),
    .Q(WX4725),
    .Q_t(WX4725_t)
  );


  nor2s3
  U2072
  (
    .DIN1(n5804),
    .DIN1_t(n5804_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX4723),
    .Q_t(WX4723_t)
  );


  nor2s3
  U2073
  (
    .DIN1(n5809),
    .DIN1_t(n5809_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX4721),
    .Q_t(WX4721_t)
  );


  nor2s3
  U2074
  (
    .DIN1(n5814),
    .DIN1_t(n5814_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX4719),
    .Q_t(WX4719_t)
  );


  nor2s3
  U2075
  (
    .DIN1(n5819),
    .DIN1_t(n5819_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX4717),
    .Q_t(WX4717_t)
  );


  nor2s3
  U2076
  (
    .DIN1(n5824),
    .DIN1_t(n5824_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX4715),
    .Q_t(WX4715_t)
  );


  nor2s3
  U2077
  (
    .DIN1(n5684),
    .DIN1_t(n5684_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX4713),
    .Q_t(WX4713_t)
  );


  nor2s3
  U2078
  (
    .DIN1(n5688),
    .DIN1_t(n5688_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX4711),
    .Q_t(WX4711_t)
  );


  nor2s3
  U2079
  (
    .DIN1(n5692),
    .DIN1_t(n5692_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX4709),
    .Q_t(WX4709_t)
  );


  nor2s3
  U2080
  (
    .DIN1(n5696),
    .DIN1_t(n5696_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX4707),
    .Q_t(WX4707_t)
  );


  nor2s3
  U2081
  (
    .DIN1(n5700),
    .DIN1_t(n5700_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX4705),
    .Q_t(WX4705_t)
  );


  nor2s3
  U2082
  (
    .DIN1(n5704),
    .DIN1_t(n5704_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX4703),
    .Q_t(WX4703_t)
  );


  nor2s3
  U2083
  (
    .DIN1(n5708),
    .DIN1_t(n5708_t),
    .DIN2(n6788),
    .DIN2_t(n6788_t),
    .Q(WX4701),
    .Q_t(WX4701_t)
  );


  nor2s3
  U2084
  (
    .DIN1(n5712),
    .DIN1_t(n5712_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX4699),
    .Q_t(WX4699_t)
  );


  nor2s3
  U2085
  (
    .DIN1(n5716),
    .DIN1_t(n5716_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX4697),
    .Q_t(WX4697_t)
  );


  nor2s3
  U2086
  (
    .DIN1(n5720),
    .DIN1_t(n5720_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX4695),
    .Q_t(WX4695_t)
  );


  nor2s3
  U2087
  (
    .DIN1(n5724),
    .DIN1_t(n5724_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX4693),
    .Q_t(WX4693_t)
  );


  nor2s3
  U2088
  (
    .DIN1(n5728),
    .DIN1_t(n5728_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX4691),
    .Q_t(WX4691_t)
  );


  nor2s3
  U2089
  (
    .DIN1(n5732),
    .DIN1_t(n5732_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX4689),
    .Q_t(WX4689_t)
  );


  nor2s3
  U2090
  (
    .DIN1(n5736),
    .DIN1_t(n5736_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX4687),
    .Q_t(WX4687_t)
  );


  nor2s3
  U2091
  (
    .DIN1(n5740),
    .DIN1_t(n5740_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX4685),
    .Q_t(WX4685_t)
  );


  nor2s3
  U2092
  (
    .DIN1(n5744),
    .DIN1_t(n5744_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX4683),
    .Q_t(WX4683_t)
  );


  and2s3
  U2093
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5748),
    .DIN2_t(n5748_t),
    .Q(WX4681),
    .Q_t(WX4681_t)
  );


  and2s3
  U2094
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5753),
    .DIN2_t(n5753_t),
    .Q(WX4679),
    .Q_t(WX4679_t)
  );


  and2s3
  U2095
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5758),
    .DIN2_t(n5758_t),
    .Q(WX4677),
    .Q_t(WX4677_t)
  );


  and2s3
  U2096
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5763),
    .DIN2_t(n5763_t),
    .Q(WX4675),
    .Q_t(WX4675_t)
  );


  and2s3
  U2097
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5768),
    .DIN2_t(n5768_t),
    .Q(WX4673),
    .Q_t(WX4673_t)
  );


  and2s3
  U2098
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5773),
    .DIN2_t(n5773_t),
    .Q(WX4671),
    .Q_t(WX4671_t)
  );


  and2s3
  U2099
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5778),
    .DIN2_t(n5778_t),
    .Q(WX4669),
    .Q_t(WX4669_t)
  );


  and2s3
  U2100
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5783),
    .DIN2_t(n5783_t),
    .Q(WX4667),
    .Q_t(WX4667_t)
  );


  and2s3
  U2101
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5788),
    .DIN2_t(n5788_t),
    .Q(WX4665),
    .Q_t(WX4665_t)
  );


  and2s3
  U2102
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5793),
    .DIN2_t(n5793_t),
    .Q(WX4663),
    .Q_t(WX4663_t)
  );


  and2s3
  U2103
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5798),
    .DIN2_t(n5798_t),
    .Q(WX4661),
    .Q_t(WX4661_t)
  );


  and2s3
  U2104
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5803),
    .DIN2_t(n5803_t),
    .Q(WX4659),
    .Q_t(WX4659_t)
  );


  and2s3
  U2105
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5808),
    .DIN2_t(n5808_t),
    .Q(WX4657),
    .Q_t(WX4657_t)
  );


  and2s3
  U2106
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5813),
    .DIN2_t(n5813_t),
    .Q(WX4655),
    .Q_t(WX4655_t)
  );


  and2s3
  U2107
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5818),
    .DIN2_t(n5818_t),
    .Q(WX4653),
    .Q_t(WX4653_t)
  );


  and2s3
  U2108
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5823),
    .DIN2_t(n5823_t),
    .Q(WX4651),
    .Q_t(WX4651_t)
  );


  and2s3
  U2109
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5683),
    .DIN2_t(n5683_t),
    .Q(WX4649),
    .Q_t(WX4649_t)
  );


  and2s3
  U2110
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5687),
    .DIN2_t(n5687_t),
    .Q(WX4647),
    .Q_t(WX4647_t)
  );


  and2s3
  U2111
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5691),
    .DIN2_t(n5691_t),
    .Q(WX4645),
    .Q_t(WX4645_t)
  );


  and2s3
  U2112
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5695),
    .DIN2_t(n5695_t),
    .Q(WX4643),
    .Q_t(WX4643_t)
  );


  and2s3
  U2113
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5699),
    .DIN2_t(n5699_t),
    .Q(WX4641),
    .Q_t(WX4641_t)
  );


  and2s3
  U2114
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5703),
    .DIN2_t(n5703_t),
    .Q(WX4639),
    .Q_t(WX4639_t)
  );


  and2s3
  U2115
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5707),
    .DIN2_t(n5707_t),
    .Q(WX4637),
    .Q_t(WX4637_t)
  );


  and2s3
  U2116
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5711),
    .DIN2_t(n5711_t),
    .Q(WX4635),
    .Q_t(WX4635_t)
  );


  and2s3
  U2117
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5715),
    .DIN2_t(n5715_t),
    .Q(WX4633),
    .Q_t(WX4633_t)
  );


  and2s3
  U2118
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5719),
    .DIN2_t(n5719_t),
    .Q(WX4631),
    .Q_t(WX4631_t)
  );


  and2s3
  U2119
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5723),
    .DIN2_t(n5723_t),
    .Q(WX4629),
    .Q_t(WX4629_t)
  );


  and2s3
  U2120
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5727),
    .DIN2_t(n5727_t),
    .Q(WX4627),
    .Q_t(WX4627_t)
  );


  and2s3
  U2121
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5731),
    .DIN2_t(n5731_t),
    .Q(WX4625),
    .Q_t(WX4625_t)
  );


  and2s3
  U2122
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5735),
    .DIN2_t(n5735_t),
    .Q(WX4623),
    .Q_t(WX4623_t)
  );


  and2s3
  U2123
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5739),
    .DIN2_t(n5739_t),
    .Q(WX4621),
    .Q_t(WX4621_t)
  );


  and2s3
  U2124
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5743),
    .DIN2_t(n5743_t),
    .Q(WX4619),
    .Q_t(WX4619_t)
  );


  nor2s3
  U2125
  (
    .DIN1(n5747),
    .DIN1_t(n5747_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX4617),
    .Q_t(WX4617_t)
  );


  nor2s3
  U2126
  (
    .DIN1(n5752),
    .DIN1_t(n5752_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX4615),
    .Q_t(WX4615_t)
  );


  nor2s3
  U2127
  (
    .DIN1(n5757),
    .DIN1_t(n5757_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX4613),
    .Q_t(WX4613_t)
  );


  nor2s3
  U2128
  (
    .DIN1(n5762),
    .DIN1_t(n5762_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX4611),
    .Q_t(WX4611_t)
  );


  nor2s3
  U2129
  (
    .DIN1(n5767),
    .DIN1_t(n5767_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4609),
    .Q_t(WX4609_t)
  );


  nor2s3
  U2130
  (
    .DIN1(n5772),
    .DIN1_t(n5772_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4607),
    .Q_t(WX4607_t)
  );


  nor2s3
  U2131
  (
    .DIN1(n5777),
    .DIN1_t(n5777_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4605),
    .Q_t(WX4605_t)
  );


  nor2s3
  U2132
  (
    .DIN1(n5782),
    .DIN1_t(n5782_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4603),
    .Q_t(WX4603_t)
  );


  nor2s3
  U2133
  (
    .DIN1(n5787),
    .DIN1_t(n5787_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4601),
    .Q_t(WX4601_t)
  );


  nor2s3
  U2134
  (
    .DIN1(n5792),
    .DIN1_t(n5792_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4599),
    .Q_t(WX4599_t)
  );


  nor2s3
  U2135
  (
    .DIN1(n5797),
    .DIN1_t(n5797_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4597),
    .Q_t(WX4597_t)
  );


  nor2s3
  U2136
  (
    .DIN1(n5802),
    .DIN1_t(n5802_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4595),
    .Q_t(WX4595_t)
  );


  nor2s3
  U2137
  (
    .DIN1(n5807),
    .DIN1_t(n5807_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4593),
    .Q_t(WX4593_t)
  );


  nor2s3
  U2138
  (
    .DIN1(n5812),
    .DIN1_t(n5812_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4591),
    .Q_t(WX4591_t)
  );


  nor2s3
  U2139
  (
    .DIN1(n5817),
    .DIN1_t(n5817_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4589),
    .Q_t(WX4589_t)
  );


  nor2s3
  U2140
  (
    .DIN1(n5822),
    .DIN1_t(n5822_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4587),
    .Q_t(WX4587_t)
  );


  nnd4s2
  U2141
  (
    .DIN1(n3684),
    .DIN1_t(n3684_t),
    .DIN2(n3685),
    .DIN2_t(n3685_t),
    .DIN3(n3686),
    .DIN3_t(n3686_t),
    .DIN4(n3687),
    .DIN4_t(n3687_t),
    .Q(WX4585),
    .Q_t(WX4585_t)
  );


  nnd2s3
  U2142
  (
    .DIN1(n3415),
    .DIN1_t(n3415_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3687),
    .Q_t(n3687_t)
  );


  xor2s3
  U2143
  (
    .DIN1(n3688),
    .DIN1_t(n3688_t),
    .DIN2(n3689),
    .DIN2_t(n3689_t),
    .Q(n3415),
    .Q_t(n3415_t)
  );


  xor2s3
  U2144
  (
    .DIN1(n5507),
    .DIN1_t(n5507_t),
    .DIN2(n5508),
    .DIN2_t(n5508_t),
    .Q(n3689),
    .Q_t(n3689_t)
  );


  xnr2s3
  U2145
  (
    .DIN1(n3253),
    .DIN1_t(n3253_t),
    .DIN2(n5509),
    .DIN2_t(n5509_t),
    .Q(n3688),
    .Q_t(n3688_t)
  );


  nnd2s3
  U2146
  (
    .DIN1(n3690),
    .DIN1_t(n3690_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3686),
    .Q_t(n3686_t)
  );


  nnd2s3
  U2147
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2081),
    .DIN2_t(n2081_t),
    .Q(n3685),
    .Q_t(n3685_t)
  );


  nnd2s3
  U2148
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n2080),
    .DIN2_t(n2080_t),
    .Q(n3684),
    .Q_t(n3684_t)
  );


  nnd4s2
  U2149
  (
    .DIN1(n3691),
    .DIN1_t(n3691_t),
    .DIN2(n3692),
    .DIN2_t(n3692_t),
    .DIN3(n3693),
    .DIN3_t(n3693_t),
    .DIN4(n3694),
    .DIN4_t(n3694_t),
    .Q(WX4583),
    .Q_t(WX4583_t)
  );


  nnd2s3
  U2150
  (
    .DIN1(n3422),
    .DIN1_t(n3422_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3694),
    .Q_t(n3694_t)
  );


  xor2s3
  U2151
  (
    .DIN1(n3695),
    .DIN1_t(n3695_t),
    .DIN2(n3696),
    .DIN2_t(n3696_t),
    .Q(n3422),
    .Q_t(n3422_t)
  );


  xor2s3
  U2152
  (
    .DIN1(n5511),
    .DIN1_t(n5511_t),
    .DIN2(n5512),
    .DIN2_t(n5512_t),
    .Q(n3696),
    .Q_t(n3696_t)
  );


  xnr2s3
  U2153
  (
    .DIN1(n3254),
    .DIN1_t(n3254_t),
    .DIN2(n5513),
    .DIN2_t(n5513_t),
    .Q(n3695),
    .Q_t(n3695_t)
  );


  nnd2s3
  U2154
  (
    .DIN1(n3697),
    .DIN1_t(n3697_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3693),
    .Q_t(n3693_t)
  );


  nnd2s3
  U2155
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2082),
    .DIN2_t(n2082_t),
    .Q(n3692),
    .Q_t(n3692_t)
  );


  nnd2s3
  U2156
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n2079),
    .DIN2_t(n2079_t),
    .Q(n3691),
    .Q_t(n3691_t)
  );


  nnd4s2
  U2157
  (
    .DIN1(n3698),
    .DIN1_t(n3698_t),
    .DIN2(n3699),
    .DIN2_t(n3699_t),
    .DIN3(n3700),
    .DIN3_t(n3700_t),
    .DIN4(n3701),
    .DIN4_t(n3701_t),
    .Q(WX4581),
    .Q_t(WX4581_t)
  );


  nnd2s3
  U2158
  (
    .DIN1(n3429),
    .DIN1_t(n3429_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3701),
    .Q_t(n3701_t)
  );


  xor2s3
  U2159
  (
    .DIN1(n3702),
    .DIN1_t(n3702_t),
    .DIN2(n3703),
    .DIN2_t(n3703_t),
    .Q(n3429),
    .Q_t(n3429_t)
  );


  xor2s3
  U2160
  (
    .DIN1(n5515),
    .DIN1_t(n5515_t),
    .DIN2(n5516),
    .DIN2_t(n5516_t),
    .Q(n3703),
    .Q_t(n3703_t)
  );


  xnr2s3
  U2161
  (
    .DIN1(n3255),
    .DIN1_t(n3255_t),
    .DIN2(n5517),
    .DIN2_t(n5517_t),
    .Q(n3702),
    .Q_t(n3702_t)
  );


  nnd2s3
  U2162
  (
    .DIN1(n3704),
    .DIN1_t(n3704_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3700),
    .Q_t(n3700_t)
  );


  nnd2s3
  U2163
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2083),
    .DIN2_t(n2083_t),
    .Q(n3699),
    .Q_t(n3699_t)
  );


  nnd2s3
  U2164
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n2078),
    .DIN2_t(n2078_t),
    .Q(n3698),
    .Q_t(n3698_t)
  );


  nnd4s2
  U2165
  (
    .DIN1(n3705),
    .DIN1_t(n3705_t),
    .DIN2(n3706),
    .DIN2_t(n3706_t),
    .DIN3(n3707),
    .DIN3_t(n3707_t),
    .DIN4(n3708),
    .DIN4_t(n3708_t),
    .Q(WX4579),
    .Q_t(WX4579_t)
  );


  nnd2s3
  U2166
  (
    .DIN1(n3436),
    .DIN1_t(n3436_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3708),
    .Q_t(n3708_t)
  );


  xor2s3
  U2167
  (
    .DIN1(n3709),
    .DIN1_t(n3709_t),
    .DIN2(n3710),
    .DIN2_t(n3710_t),
    .Q(n3436),
    .Q_t(n3436_t)
  );


  xor2s3
  U2168
  (
    .DIN1(n5519),
    .DIN1_t(n5519_t),
    .DIN2(n5520),
    .DIN2_t(n5520_t),
    .Q(n3710),
    .Q_t(n3710_t)
  );


  xnr2s3
  U2169
  (
    .DIN1(n3256),
    .DIN1_t(n3256_t),
    .DIN2(n5521),
    .DIN2_t(n5521_t),
    .Q(n3709),
    .Q_t(n3709_t)
  );


  nnd2s3
  U2170
  (
    .DIN1(n3711),
    .DIN1_t(n3711_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3707),
    .Q_t(n3707_t)
  );


  nnd2s3
  U2171
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2084),
    .DIN2_t(n2084_t),
    .Q(n3706),
    .Q_t(n3706_t)
  );


  nnd2s3
  U2172
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n2077),
    .DIN2_t(n2077_t),
    .Q(n3705),
    .Q_t(n3705_t)
  );


  nnd4s2
  U2173
  (
    .DIN1(n3712),
    .DIN1_t(n3712_t),
    .DIN2(n3713),
    .DIN2_t(n3713_t),
    .DIN3(n3714),
    .DIN3_t(n3714_t),
    .DIN4(n3715),
    .DIN4_t(n3715_t),
    .Q(WX4577),
    .Q_t(WX4577_t)
  );


  nnd2s3
  U2174
  (
    .DIN1(n3443),
    .DIN1_t(n3443_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3715),
    .Q_t(n3715_t)
  );


  xor2s3
  U2175
  (
    .DIN1(n3716),
    .DIN1_t(n3716_t),
    .DIN2(n3717),
    .DIN2_t(n3717_t),
    .Q(n3443),
    .Q_t(n3443_t)
  );


  xor2s3
  U2176
  (
    .DIN1(n5523),
    .DIN1_t(n5523_t),
    .DIN2(n5524),
    .DIN2_t(n5524_t),
    .Q(n3717),
    .Q_t(n3717_t)
  );


  xnr2s3
  U2177
  (
    .DIN1(n3257),
    .DIN1_t(n3257_t),
    .DIN2(n5525),
    .DIN2_t(n5525_t),
    .Q(n3716),
    .Q_t(n3716_t)
  );


  nnd2s3
  U2178
  (
    .DIN1(n3718),
    .DIN1_t(n3718_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3714),
    .Q_t(n3714_t)
  );


  nnd2s3
  U2179
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2085),
    .DIN2_t(n2085_t),
    .Q(n3713),
    .Q_t(n3713_t)
  );


  nnd2s3
  U2180
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n2076),
    .DIN2_t(n2076_t),
    .Q(n3712),
    .Q_t(n3712_t)
  );


  nnd4s2
  U2181
  (
    .DIN1(n3719),
    .DIN1_t(n3719_t),
    .DIN2(n3720),
    .DIN2_t(n3720_t),
    .DIN3(n3721),
    .DIN3_t(n3721_t),
    .DIN4(n3722),
    .DIN4_t(n3722_t),
    .Q(WX4575),
    .Q_t(WX4575_t)
  );


  nnd2s3
  U2182
  (
    .DIN1(n3450),
    .DIN1_t(n3450_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3722),
    .Q_t(n3722_t)
  );


  xor2s3
  U2183
  (
    .DIN1(n3723),
    .DIN1_t(n3723_t),
    .DIN2(n3724),
    .DIN2_t(n3724_t),
    .Q(n3450),
    .Q_t(n3450_t)
  );


  xor2s3
  U2184
  (
    .DIN1(n5527),
    .DIN1_t(n5527_t),
    .DIN2(n5528),
    .DIN2_t(n5528_t),
    .Q(n3724),
    .Q_t(n3724_t)
  );


  xnr2s3
  U2185
  (
    .DIN1(n3258),
    .DIN1_t(n3258_t),
    .DIN2(n5529),
    .DIN2_t(n5529_t),
    .Q(n3723),
    .Q_t(n3723_t)
  );


  nnd2s3
  U2186
  (
    .DIN1(n3725),
    .DIN1_t(n3725_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3721),
    .Q_t(n3721_t)
  );


  nnd2s3
  U2187
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2086),
    .DIN2_t(n2086_t),
    .Q(n3720),
    .Q_t(n3720_t)
  );


  nnd2s3
  U2188
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n2075),
    .DIN2_t(n2075_t),
    .Q(n3719),
    .Q_t(n3719_t)
  );


  nnd4s2
  U2189
  (
    .DIN1(n3726),
    .DIN1_t(n3726_t),
    .DIN2(n3727),
    .DIN2_t(n3727_t),
    .DIN3(n3728),
    .DIN3_t(n3728_t),
    .DIN4(n3729),
    .DIN4_t(n3729_t),
    .Q(WX4573),
    .Q_t(WX4573_t)
  );


  nnd2s3
  U2190
  (
    .DIN1(n3457),
    .DIN1_t(n3457_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3729),
    .Q_t(n3729_t)
  );


  xor2s3
  U2191
  (
    .DIN1(n3730),
    .DIN1_t(n3730_t),
    .DIN2(n3731),
    .DIN2_t(n3731_t),
    .Q(n3457),
    .Q_t(n3457_t)
  );


  xor2s3
  U2192
  (
    .DIN1(n5531),
    .DIN1_t(n5531_t),
    .DIN2(n5532),
    .DIN2_t(n5532_t),
    .Q(n3731),
    .Q_t(n3731_t)
  );


  xnr2s3
  U2193
  (
    .DIN1(n3259),
    .DIN1_t(n3259_t),
    .DIN2(n5533),
    .DIN2_t(n5533_t),
    .Q(n3730),
    .Q_t(n3730_t)
  );


  nnd2s3
  U2194
  (
    .DIN1(n3732),
    .DIN1_t(n3732_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3728),
    .Q_t(n3728_t)
  );


  nnd2s3
  U2195
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2087),
    .DIN2_t(n2087_t),
    .Q(n3727),
    .Q_t(n3727_t)
  );


  nnd2s3
  U2196
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n2074),
    .DIN2_t(n2074_t),
    .Q(n3726),
    .Q_t(n3726_t)
  );


  nnd4s2
  U2197
  (
    .DIN1(n3733),
    .DIN1_t(n3733_t),
    .DIN2(n3734),
    .DIN2_t(n3734_t),
    .DIN3(n3735),
    .DIN3_t(n3735_t),
    .DIN4(n3736),
    .DIN4_t(n3736_t),
    .Q(WX4571),
    .Q_t(WX4571_t)
  );


  nnd2s3
  U2198
  (
    .DIN1(n3464),
    .DIN1_t(n3464_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3736),
    .Q_t(n3736_t)
  );


  xor2s3
  U2199
  (
    .DIN1(n3737),
    .DIN1_t(n3737_t),
    .DIN2(n3738),
    .DIN2_t(n3738_t),
    .Q(n3464),
    .Q_t(n3464_t)
  );


  xor2s3
  U2200
  (
    .DIN1(n5535),
    .DIN1_t(n5535_t),
    .DIN2(n5536),
    .DIN2_t(n5536_t),
    .Q(n3738),
    .Q_t(n3738_t)
  );


  xnr2s3
  U2201
  (
    .DIN1(n3260),
    .DIN1_t(n3260_t),
    .DIN2(n5537),
    .DIN2_t(n5537_t),
    .Q(n3737),
    .Q_t(n3737_t)
  );


  nnd2s3
  U2202
  (
    .DIN1(n3739),
    .DIN1_t(n3739_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3735),
    .Q_t(n3735_t)
  );


  nnd2s3
  U2203
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2088),
    .DIN2_t(n2088_t),
    .Q(n3734),
    .Q_t(n3734_t)
  );


  nnd2s3
  U2204
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n2073),
    .DIN2_t(n2073_t),
    .Q(n3733),
    .Q_t(n3733_t)
  );


  nnd4s2
  U2205
  (
    .DIN1(n3740),
    .DIN1_t(n3740_t),
    .DIN2(n3741),
    .DIN2_t(n3741_t),
    .DIN3(n3742),
    .DIN3_t(n3742_t),
    .DIN4(n3743),
    .DIN4_t(n3743_t),
    .Q(WX4569),
    .Q_t(WX4569_t)
  );


  nnd2s3
  U2206
  (
    .DIN1(n3471),
    .DIN1_t(n3471_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3743),
    .Q_t(n3743_t)
  );


  xor2s3
  U2207
  (
    .DIN1(n3744),
    .DIN1_t(n3744_t),
    .DIN2(n3745),
    .DIN2_t(n3745_t),
    .Q(n3471),
    .Q_t(n3471_t)
  );


  xor2s3
  U2208
  (
    .DIN1(n5539),
    .DIN1_t(n5539_t),
    .DIN2(n5540),
    .DIN2_t(n5540_t),
    .Q(n3745),
    .Q_t(n3745_t)
  );


  xnr2s3
  U2209
  (
    .DIN1(n3261),
    .DIN1_t(n3261_t),
    .DIN2(n5541),
    .DIN2_t(n5541_t),
    .Q(n3744),
    .Q_t(n3744_t)
  );


  nnd2s3
  U2210
  (
    .DIN1(n3746),
    .DIN1_t(n3746_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3742),
    .Q_t(n3742_t)
  );


  nnd2s3
  U2211
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2089),
    .DIN2_t(n2089_t),
    .Q(n3741),
    .Q_t(n3741_t)
  );


  nnd2s3
  U2212
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n2072),
    .DIN2_t(n2072_t),
    .Q(n3740),
    .Q_t(n3740_t)
  );


  nnd4s2
  U2213
  (
    .DIN1(n3747),
    .DIN1_t(n3747_t),
    .DIN2(n3748),
    .DIN2_t(n3748_t),
    .DIN3(n3749),
    .DIN3_t(n3749_t),
    .DIN4(n3750),
    .DIN4_t(n3750_t),
    .Q(WX4567),
    .Q_t(WX4567_t)
  );


  nnd2s3
  U2214
  (
    .DIN1(n3478),
    .DIN1_t(n3478_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3750),
    .Q_t(n3750_t)
  );


  xor2s3
  U2215
  (
    .DIN1(n3751),
    .DIN1_t(n3751_t),
    .DIN2(n3752),
    .DIN2_t(n3752_t),
    .Q(n3478),
    .Q_t(n3478_t)
  );


  xor2s3
  U2216
  (
    .DIN1(n5543),
    .DIN1_t(n5543_t),
    .DIN2(n5544),
    .DIN2_t(n5544_t),
    .Q(n3752),
    .Q_t(n3752_t)
  );


  xnr2s3
  U2217
  (
    .DIN1(n3262),
    .DIN1_t(n3262_t),
    .DIN2(n5545),
    .DIN2_t(n5545_t),
    .Q(n3751),
    .Q_t(n3751_t)
  );


  nnd2s3
  U2218
  (
    .DIN1(n3753),
    .DIN1_t(n3753_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3749),
    .Q_t(n3749_t)
  );


  nnd2s3
  U2219
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2090),
    .DIN2_t(n2090_t),
    .Q(n3748),
    .Q_t(n3748_t)
  );


  nnd2s3
  U2220
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n2071),
    .DIN2_t(n2071_t),
    .Q(n3747),
    .Q_t(n3747_t)
  );


  nnd4s2
  U2221
  (
    .DIN1(n3754),
    .DIN1_t(n3754_t),
    .DIN2(n3755),
    .DIN2_t(n3755_t),
    .DIN3(n3756),
    .DIN3_t(n3756_t),
    .DIN4(n3757),
    .DIN4_t(n3757_t),
    .Q(WX4565),
    .Q_t(WX4565_t)
  );


  nnd2s3
  U2222
  (
    .DIN1(n3485),
    .DIN1_t(n3485_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3757),
    .Q_t(n3757_t)
  );


  xor2s3
  U2223
  (
    .DIN1(n3758),
    .DIN1_t(n3758_t),
    .DIN2(n3759),
    .DIN2_t(n3759_t),
    .Q(n3485),
    .Q_t(n3485_t)
  );


  xor2s3
  U2224
  (
    .DIN1(n5547),
    .DIN1_t(n5547_t),
    .DIN2(n5548),
    .DIN2_t(n5548_t),
    .Q(n3759),
    .Q_t(n3759_t)
  );


  xnr2s3
  U2225
  (
    .DIN1(n3263),
    .DIN1_t(n3263_t),
    .DIN2(n5549),
    .DIN2_t(n5549_t),
    .Q(n3758),
    .Q_t(n3758_t)
  );


  nnd2s3
  U2226
  (
    .DIN1(n3760),
    .DIN1_t(n3760_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3756),
    .Q_t(n3756_t)
  );


  nnd2s3
  U2227
  (
    .DIN1(n6603),
    .DIN1_t(n6603_t),
    .DIN2(n2091),
    .DIN2_t(n2091_t),
    .Q(n3755),
    .Q_t(n3755_t)
  );


  nnd2s3
  U2228
  (
    .DIN1(n6572),
    .DIN1_t(n6572_t),
    .DIN2(n2070),
    .DIN2_t(n2070_t),
    .Q(n3754),
    .Q_t(n3754_t)
  );


  nnd4s2
  U2229
  (
    .DIN1(n3761),
    .DIN1_t(n3761_t),
    .DIN2(n3762),
    .DIN2_t(n3762_t),
    .DIN3(n3763),
    .DIN3_t(n3763_t),
    .DIN4(n3764),
    .DIN4_t(n3764_t),
    .Q(WX4563),
    .Q_t(WX4563_t)
  );


  nnd2s3
  U2230
  (
    .DIN1(n3492),
    .DIN1_t(n3492_t),
    .DIN2(n6645),
    .DIN2_t(n6645_t),
    .Q(n3764),
    .Q_t(n3764_t)
  );


  xor2s3
  U2231
  (
    .DIN1(n3765),
    .DIN1_t(n3765_t),
    .DIN2(n3766),
    .DIN2_t(n3766_t),
    .Q(n3492),
    .Q_t(n3492_t)
  );


  xor2s3
  U2232
  (
    .DIN1(n5551),
    .DIN1_t(n5551_t),
    .DIN2(n5552),
    .DIN2_t(n5552_t),
    .Q(n3766),
    .Q_t(n3766_t)
  );


  xnr2s3
  U2233
  (
    .DIN1(n3264),
    .DIN1_t(n3264_t),
    .DIN2(n5553),
    .DIN2_t(n5553_t),
    .Q(n3765),
    .Q_t(n3765_t)
  );


  nnd2s3
  U2234
  (
    .DIN1(n3767),
    .DIN1_t(n3767_t),
    .DIN2(n6676),
    .DIN2_t(n6676_t),
    .Q(n3763),
    .Q_t(n3763_t)
  );


  nnd2s3
  U2235
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2092),
    .DIN2_t(n2092_t),
    .Q(n3762),
    .Q_t(n3762_t)
  );


  nnd2s3
  U2236
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2069),
    .DIN2_t(n2069_t),
    .Q(n3761),
    .Q_t(n3761_t)
  );


  nnd4s2
  U2237
  (
    .DIN1(n3768),
    .DIN1_t(n3768_t),
    .DIN2(n3769),
    .DIN2_t(n3769_t),
    .DIN3(n3770),
    .DIN3_t(n3770_t),
    .DIN4(n3771),
    .DIN4_t(n3771_t),
    .Q(WX4561),
    .Q_t(WX4561_t)
  );


  nnd2s3
  U2238
  (
    .DIN1(n3499),
    .DIN1_t(n3499_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3771),
    .Q_t(n3771_t)
  );


  xor2s3
  U2239
  (
    .DIN1(n3772),
    .DIN1_t(n3772_t),
    .DIN2(n3773),
    .DIN2_t(n3773_t),
    .Q(n3499),
    .Q_t(n3499_t)
  );


  xor2s3
  U2240
  (
    .DIN1(n5555),
    .DIN1_t(n5555_t),
    .DIN2(n5556),
    .DIN2_t(n5556_t),
    .Q(n3773),
    .Q_t(n3773_t)
  );


  xnr2s3
  U2241
  (
    .DIN1(n3265),
    .DIN1_t(n3265_t),
    .DIN2(n5557),
    .DIN2_t(n5557_t),
    .Q(n3772),
    .Q_t(n3772_t)
  );


  nnd2s3
  U2242
  (
    .DIN1(n3774),
    .DIN1_t(n3774_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3770),
    .Q_t(n3770_t)
  );


  nnd2s3
  U2243
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2093),
    .DIN2_t(n2093_t),
    .Q(n3769),
    .Q_t(n3769_t)
  );


  nnd2s3
  U2244
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2068),
    .DIN2_t(n2068_t),
    .Q(n3768),
    .Q_t(n3768_t)
  );


  nnd4s2
  U2245
  (
    .DIN1(n3775),
    .DIN1_t(n3775_t),
    .DIN2(n3776),
    .DIN2_t(n3776_t),
    .DIN3(n3777),
    .DIN3_t(n3777_t),
    .DIN4(n3778),
    .DIN4_t(n3778_t),
    .Q(WX4559),
    .Q_t(WX4559_t)
  );


  nnd2s3
  U2246
  (
    .DIN1(n3506),
    .DIN1_t(n3506_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3778),
    .Q_t(n3778_t)
  );


  xor2s3
  U2247
  (
    .DIN1(n3779),
    .DIN1_t(n3779_t),
    .DIN2(n3780),
    .DIN2_t(n3780_t),
    .Q(n3506),
    .Q_t(n3506_t)
  );


  xor2s3
  U2248
  (
    .DIN1(n5559),
    .DIN1_t(n5559_t),
    .DIN2(n5560),
    .DIN2_t(n5560_t),
    .Q(n3780),
    .Q_t(n3780_t)
  );


  xnr2s3
  U2249
  (
    .DIN1(n3266),
    .DIN1_t(n3266_t),
    .DIN2(n5561),
    .DIN2_t(n5561_t),
    .Q(n3779),
    .Q_t(n3779_t)
  );


  nnd2s3
  U2250
  (
    .DIN1(n3781),
    .DIN1_t(n3781_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3777),
    .Q_t(n3777_t)
  );


  nnd2s3
  U2251
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2094),
    .DIN2_t(n2094_t),
    .Q(n3776),
    .Q_t(n3776_t)
  );


  nnd2s3
  U2252
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2067),
    .DIN2_t(n2067_t),
    .Q(n3775),
    .Q_t(n3775_t)
  );


  nnd4s2
  U2253
  (
    .DIN1(n3782),
    .DIN1_t(n3782_t),
    .DIN2(n3783),
    .DIN2_t(n3783_t),
    .DIN3(n3784),
    .DIN3_t(n3784_t),
    .DIN4(n3785),
    .DIN4_t(n3785_t),
    .Q(WX4557),
    .Q_t(WX4557_t)
  );


  nnd2s3
  U2254
  (
    .DIN1(n3513),
    .DIN1_t(n3513_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3785),
    .Q_t(n3785_t)
  );


  xor2s3
  U2255
  (
    .DIN1(n3786),
    .DIN1_t(n3786_t),
    .DIN2(n3787),
    .DIN2_t(n3787_t),
    .Q(n3513),
    .Q_t(n3513_t)
  );


  xor2s3
  U2256
  (
    .DIN1(n5563),
    .DIN1_t(n5563_t),
    .DIN2(n5564),
    .DIN2_t(n5564_t),
    .Q(n3787),
    .Q_t(n3787_t)
  );


  xnr2s3
  U2257
  (
    .DIN1(n3267),
    .DIN1_t(n3267_t),
    .DIN2(n5565),
    .DIN2_t(n5565_t),
    .Q(n3786),
    .Q_t(n3786_t)
  );


  nnd2s3
  U2258
  (
    .DIN1(n3788),
    .DIN1_t(n3788_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3784),
    .Q_t(n3784_t)
  );


  nnd2s3
  U2259
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2095),
    .DIN2_t(n2095_t),
    .Q(n3783),
    .Q_t(n3783_t)
  );


  nnd2s3
  U2260
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2066),
    .DIN2_t(n2066_t),
    .Q(n3782),
    .Q_t(n3782_t)
  );


  nnd4s2
  U2261
  (
    .DIN1(n3789),
    .DIN1_t(n3789_t),
    .DIN2(n3790),
    .DIN2_t(n3790_t),
    .DIN3(n3791),
    .DIN3_t(n3791_t),
    .DIN4(n3792),
    .DIN4_t(n3792_t),
    .Q(WX4555),
    .Q_t(WX4555_t)
  );


  nnd2s3
  U2262
  (
    .DIN1(n3520),
    .DIN1_t(n3520_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3792),
    .Q_t(n3792_t)
  );


  xor2s3
  U2263
  (
    .DIN1(n3793),
    .DIN1_t(n3793_t),
    .DIN2(n3794),
    .DIN2_t(n3794_t),
    .Q(n3520),
    .Q_t(n3520_t)
  );


  xor2s3
  U2264
  (
    .DIN1(n5567),
    .DIN1_t(n5567_t),
    .DIN2(n5568),
    .DIN2_t(n5568_t),
    .Q(n3794),
    .Q_t(n3794_t)
  );


  xnr2s3
  U2265
  (
    .DIN1(n3268),
    .DIN1_t(n3268_t),
    .DIN2(n5569),
    .DIN2_t(n5569_t),
    .Q(n3793),
    .Q_t(n3793_t)
  );


  nnd2s3
  U2266
  (
    .DIN1(n3795),
    .DIN1_t(n3795_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3791),
    .Q_t(n3791_t)
  );


  nnd2s3
  U2267
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2096),
    .DIN2_t(n2096_t),
    .Q(n3790),
    .Q_t(n3790_t)
  );


  nnd2s3
  U2268
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2065),
    .DIN2_t(n2065_t),
    .Q(n3789),
    .Q_t(n3789_t)
  );


  nnd4s2
  U2269
  (
    .DIN1(n3796),
    .DIN1_t(n3796_t),
    .DIN2(n3797),
    .DIN2_t(n3797_t),
    .DIN3(n3798),
    .DIN3_t(n3798_t),
    .DIN4(n3799),
    .DIN4_t(n3799_t),
    .Q(WX4553),
    .Q_t(WX4553_t)
  );


  nnd2s3
  U2270
  (
    .DIN1(n3528),
    .DIN1_t(n3528_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3799),
    .Q_t(n3799_t)
  );


  xor2s3
  U2271
  (
    .DIN1(n3800),
    .DIN1_t(n3800_t),
    .DIN2(n3801),
    .DIN2_t(n3801_t),
    .Q(n3528),
    .Q_t(n3528_t)
  );


  xor2s3
  U2272
  (
    .DIN1(n5573),
    .DIN1_t(n5573_t),
    .DIN2(n3802),
    .DIN2_t(n3802_t),
    .Q(n3801),
    .Q_t(n3801_t)
  );


  xor2s3
  U2273
  (
    .DIN1(n5571),
    .DIN1_t(n5571_t),
    .DIN2(n5572),
    .DIN2_t(n5572_t),
    .Q(n3802),
    .Q_t(n3802_t)
  );


  xor2s3
  U2274
  (
    .DIN1(n5574),
    .DIN1_t(n5574_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3800),
    .Q_t(n3800_t)
  );


  nnd2s3
  U2275
  (
    .DIN1(n3803),
    .DIN1_t(n3803_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3798),
    .Q_t(n3798_t)
  );


  nnd2s3
  U2276
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2097),
    .DIN2_t(n2097_t),
    .Q(n3797),
    .Q_t(n3797_t)
  );


  nnd2s3
  U2277
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2064),
    .DIN2_t(n2064_t),
    .Q(n3796),
    .Q_t(n3796_t)
  );


  nnd4s2
  U2278
  (
    .DIN1(n3804),
    .DIN1_t(n3804_t),
    .DIN2(n3805),
    .DIN2_t(n3805_t),
    .DIN3(n3806),
    .DIN3_t(n3806_t),
    .DIN4(n3807),
    .DIN4_t(n3807_t),
    .Q(WX4551),
    .Q_t(WX4551_t)
  );


  nnd2s3
  U2279
  (
    .DIN1(n3536),
    .DIN1_t(n3536_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3807),
    .Q_t(n3807_t)
  );


  xor2s3
  U2280
  (
    .DIN1(n3808),
    .DIN1_t(n3808_t),
    .DIN2(n3809),
    .DIN2_t(n3809_t),
    .Q(n3536),
    .Q_t(n3536_t)
  );


  xor2s3
  U2281
  (
    .DIN1(n5578),
    .DIN1_t(n5578_t),
    .DIN2(n3810),
    .DIN2_t(n3810_t),
    .Q(n3809),
    .Q_t(n3809_t)
  );


  xor2s3
  U2282
  (
    .DIN1(n5576),
    .DIN1_t(n5576_t),
    .DIN2(n5577),
    .DIN2_t(n5577_t),
    .Q(n3810),
    .Q_t(n3810_t)
  );


  xor2s3
  U2283
  (
    .DIN1(n5579),
    .DIN1_t(n5579_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3808),
    .Q_t(n3808_t)
  );


  nnd2s3
  U2284
  (
    .DIN1(n3811),
    .DIN1_t(n3811_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3806),
    .Q_t(n3806_t)
  );


  nnd2s3
  U2285
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2098),
    .DIN2_t(n2098_t),
    .Q(n3805),
    .Q_t(n3805_t)
  );


  nnd2s3
  U2286
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2063),
    .DIN2_t(n2063_t),
    .Q(n3804),
    .Q_t(n3804_t)
  );


  nnd4s2
  U2287
  (
    .DIN1(n3812),
    .DIN1_t(n3812_t),
    .DIN2(n3813),
    .DIN2_t(n3813_t),
    .DIN3(n3814),
    .DIN3_t(n3814_t),
    .DIN4(n3815),
    .DIN4_t(n3815_t),
    .Q(WX4549),
    .Q_t(WX4549_t)
  );


  nnd2s3
  U2288
  (
    .DIN1(n3544),
    .DIN1_t(n3544_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3815),
    .Q_t(n3815_t)
  );


  xor2s3
  U2289
  (
    .DIN1(n3816),
    .DIN1_t(n3816_t),
    .DIN2(n3817),
    .DIN2_t(n3817_t),
    .Q(n3544),
    .Q_t(n3544_t)
  );


  xor2s3
  U2290
  (
    .DIN1(n5583),
    .DIN1_t(n5583_t),
    .DIN2(n3818),
    .DIN2_t(n3818_t),
    .Q(n3817),
    .Q_t(n3817_t)
  );


  xor2s3
  U2291
  (
    .DIN1(n5581),
    .DIN1_t(n5581_t),
    .DIN2(n5582),
    .DIN2_t(n5582_t),
    .Q(n3818),
    .Q_t(n3818_t)
  );


  xor2s3
  U2292
  (
    .DIN1(n5584),
    .DIN1_t(n5584_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3816),
    .Q_t(n3816_t)
  );


  nnd2s3
  U2293
  (
    .DIN1(n3819),
    .DIN1_t(n3819_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3814),
    .Q_t(n3814_t)
  );


  nnd2s3
  U2294
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2099),
    .DIN2_t(n2099_t),
    .Q(n3813),
    .Q_t(n3813_t)
  );


  nnd2s3
  U2295
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2062),
    .DIN2_t(n2062_t),
    .Q(n3812),
    .Q_t(n3812_t)
  );


  nnd4s2
  U2296
  (
    .DIN1(n3820),
    .DIN1_t(n3820_t),
    .DIN2(n3821),
    .DIN2_t(n3821_t),
    .DIN3(n3822),
    .DIN3_t(n3822_t),
    .DIN4(n3823),
    .DIN4_t(n3823_t),
    .Q(WX4547),
    .Q_t(WX4547_t)
  );


  nnd2s3
  U2297
  (
    .DIN1(n3552),
    .DIN1_t(n3552_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3823),
    .Q_t(n3823_t)
  );


  xor2s3
  U2298
  (
    .DIN1(n3824),
    .DIN1_t(n3824_t),
    .DIN2(n3825),
    .DIN2_t(n3825_t),
    .Q(n3552),
    .Q_t(n3552_t)
  );


  xor2s3
  U2299
  (
    .DIN1(n5588),
    .DIN1_t(n5588_t),
    .DIN2(n3826),
    .DIN2_t(n3826_t),
    .Q(n3825),
    .Q_t(n3825_t)
  );


  xor2s3
  U2300
  (
    .DIN1(n5586),
    .DIN1_t(n5586_t),
    .DIN2(n5587),
    .DIN2_t(n5587_t),
    .Q(n3826),
    .Q_t(n3826_t)
  );


  xor2s3
  U2301
  (
    .DIN1(n5589),
    .DIN1_t(n5589_t),
    .DIN2(n6690),
    .DIN2_t(n6690_t),
    .Q(n3824),
    .Q_t(n3824_t)
  );


  nnd2s3
  U2302
  (
    .DIN1(n3827),
    .DIN1_t(n3827_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3822),
    .Q_t(n3822_t)
  );


  nnd2s3
  U2303
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2100),
    .DIN2_t(n2100_t),
    .Q(n3821),
    .Q_t(n3821_t)
  );


  nnd2s3
  U2304
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2061),
    .DIN2_t(n2061_t),
    .Q(n3820),
    .Q_t(n3820_t)
  );


  nnd4s2
  U2305
  (
    .DIN1(n3828),
    .DIN1_t(n3828_t),
    .DIN2(n3829),
    .DIN2_t(n3829_t),
    .DIN3(n3830),
    .DIN3_t(n3830_t),
    .DIN4(n3831),
    .DIN4_t(n3831_t),
    .Q(WX4545),
    .Q_t(WX4545_t)
  );


  nnd2s3
  U2306
  (
    .DIN1(n3560),
    .DIN1_t(n3560_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3831),
    .Q_t(n3831_t)
  );


  xor2s3
  U2307
  (
    .DIN1(n3832),
    .DIN1_t(n3832_t),
    .DIN2(n3833),
    .DIN2_t(n3833_t),
    .Q(n3560),
    .Q_t(n3560_t)
  );


  xor2s3
  U2308
  (
    .DIN1(n5593),
    .DIN1_t(n5593_t),
    .DIN2(n3834),
    .DIN2_t(n3834_t),
    .Q(n3833),
    .Q_t(n3833_t)
  );


  xor2s3
  U2309
  (
    .DIN1(n5591),
    .DIN1_t(n5591_t),
    .DIN2(n5592),
    .DIN2_t(n5592_t),
    .Q(n3834),
    .Q_t(n3834_t)
  );


  xor2s3
  U2310
  (
    .DIN1(n5594),
    .DIN1_t(n5594_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3832),
    .Q_t(n3832_t)
  );


  nnd2s3
  U2311
  (
    .DIN1(n3835),
    .DIN1_t(n3835_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3830),
    .Q_t(n3830_t)
  );


  nnd2s3
  U2312
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2101),
    .DIN2_t(n2101_t),
    .Q(n3829),
    .Q_t(n3829_t)
  );


  nnd2s3
  U2313
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2060),
    .DIN2_t(n2060_t),
    .Q(n3828),
    .Q_t(n3828_t)
  );


  nnd4s2
  U2314
  (
    .DIN1(n3836),
    .DIN1_t(n3836_t),
    .DIN2(n3837),
    .DIN2_t(n3837_t),
    .DIN3(n3838),
    .DIN3_t(n3838_t),
    .DIN4(n3839),
    .DIN4_t(n3839_t),
    .Q(WX4543),
    .Q_t(WX4543_t)
  );


  nnd2s3
  U2315
  (
    .DIN1(n3568),
    .DIN1_t(n3568_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3839),
    .Q_t(n3839_t)
  );


  xor2s3
  U2316
  (
    .DIN1(n3840),
    .DIN1_t(n3840_t),
    .DIN2(n3841),
    .DIN2_t(n3841_t),
    .Q(n3568),
    .Q_t(n3568_t)
  );


  xor2s3
  U2317
  (
    .DIN1(n5598),
    .DIN1_t(n5598_t),
    .DIN2(n3842),
    .DIN2_t(n3842_t),
    .Q(n3841),
    .Q_t(n3841_t)
  );


  xor2s3
  U2318
  (
    .DIN1(n5596),
    .DIN1_t(n5596_t),
    .DIN2(n5597),
    .DIN2_t(n5597_t),
    .Q(n3842),
    .Q_t(n3842_t)
  );


  xor2s3
  U2319
  (
    .DIN1(n5599),
    .DIN1_t(n5599_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3840),
    .Q_t(n3840_t)
  );


  nnd2s3
  U2320
  (
    .DIN1(n3843),
    .DIN1_t(n3843_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3838),
    .Q_t(n3838_t)
  );


  nnd2s3
  U2321
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2102),
    .DIN2_t(n2102_t),
    .Q(n3837),
    .Q_t(n3837_t)
  );


  nnd2s3
  U2322
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2059),
    .DIN2_t(n2059_t),
    .Q(n3836),
    .Q_t(n3836_t)
  );


  nnd4s2
  U2323
  (
    .DIN1(n3844),
    .DIN1_t(n3844_t),
    .DIN2(n3845),
    .DIN2_t(n3845_t),
    .DIN3(n3846),
    .DIN3_t(n3846_t),
    .DIN4(n3847),
    .DIN4_t(n3847_t),
    .Q(WX4541),
    .Q_t(WX4541_t)
  );


  nnd2s3
  U2324
  (
    .DIN1(n3576),
    .DIN1_t(n3576_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3847),
    .Q_t(n3847_t)
  );


  xor2s3
  U2325
  (
    .DIN1(n3848),
    .DIN1_t(n3848_t),
    .DIN2(n3849),
    .DIN2_t(n3849_t),
    .Q(n3576),
    .Q_t(n3576_t)
  );


  xor2s3
  U2326
  (
    .DIN1(n5603),
    .DIN1_t(n5603_t),
    .DIN2(n3850),
    .DIN2_t(n3850_t),
    .Q(n3849),
    .Q_t(n3849_t)
  );


  xor2s3
  U2327
  (
    .DIN1(n5601),
    .DIN1_t(n5601_t),
    .DIN2(n5602),
    .DIN2_t(n5602_t),
    .Q(n3850),
    .Q_t(n3850_t)
  );


  xor2s3
  U2328
  (
    .DIN1(n5604),
    .DIN1_t(n5604_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3848),
    .Q_t(n3848_t)
  );


  nnd2s3
  U2329
  (
    .DIN1(n3851),
    .DIN1_t(n3851_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3846),
    .Q_t(n3846_t)
  );


  nnd2s3
  U2330
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2103),
    .DIN2_t(n2103_t),
    .Q(n3845),
    .Q_t(n3845_t)
  );


  nnd2s3
  U2331
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2058),
    .DIN2_t(n2058_t),
    .Q(n3844),
    .Q_t(n3844_t)
  );


  nnd4s2
  U2332
  (
    .DIN1(n3852),
    .DIN1_t(n3852_t),
    .DIN2(n3853),
    .DIN2_t(n3853_t),
    .DIN3(n3854),
    .DIN3_t(n3854_t),
    .DIN4(n3855),
    .DIN4_t(n3855_t),
    .Q(WX4539),
    .Q_t(WX4539_t)
  );


  nnd2s3
  U2333
  (
    .DIN1(n3584),
    .DIN1_t(n3584_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3855),
    .Q_t(n3855_t)
  );


  xor2s3
  U2334
  (
    .DIN1(n3856),
    .DIN1_t(n3856_t),
    .DIN2(n3857),
    .DIN2_t(n3857_t),
    .Q(n3584),
    .Q_t(n3584_t)
  );


  xor2s3
  U2335
  (
    .DIN1(n5608),
    .DIN1_t(n5608_t),
    .DIN2(n3858),
    .DIN2_t(n3858_t),
    .Q(n3857),
    .Q_t(n3857_t)
  );


  xor2s3
  U2336
  (
    .DIN1(n5606),
    .DIN1_t(n5606_t),
    .DIN2(n5607),
    .DIN2_t(n5607_t),
    .Q(n3858),
    .Q_t(n3858_t)
  );


  xor2s3
  U2337
  (
    .DIN1(n5609),
    .DIN1_t(n5609_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3856),
    .Q_t(n3856_t)
  );


  nnd2s3
  U2338
  (
    .DIN1(n3859),
    .DIN1_t(n3859_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3854),
    .Q_t(n3854_t)
  );


  nnd2s3
  U2339
  (
    .DIN1(n6602),
    .DIN1_t(n6602_t),
    .DIN2(n2104),
    .DIN2_t(n2104_t),
    .Q(n3853),
    .Q_t(n3853_t)
  );


  nnd2s3
  U2340
  (
    .DIN1(n6571),
    .DIN1_t(n6571_t),
    .DIN2(n2057),
    .DIN2_t(n2057_t),
    .Q(n3852),
    .Q_t(n3852_t)
  );


  nnd4s2
  U2341
  (
    .DIN1(n3860),
    .DIN1_t(n3860_t),
    .DIN2(n3861),
    .DIN2_t(n3861_t),
    .DIN3(n3862),
    .DIN3_t(n3862_t),
    .DIN4(n3863),
    .DIN4_t(n3863_t),
    .Q(WX4537),
    .Q_t(WX4537_t)
  );


  nnd2s3
  U2342
  (
    .DIN1(n3592),
    .DIN1_t(n3592_t),
    .DIN2(n6644),
    .DIN2_t(n6644_t),
    .Q(n3863),
    .Q_t(n3863_t)
  );


  xor2s3
  U2343
  (
    .DIN1(n3864),
    .DIN1_t(n3864_t),
    .DIN2(n3865),
    .DIN2_t(n3865_t),
    .Q(n3592),
    .Q_t(n3592_t)
  );


  xor2s3
  U2344
  (
    .DIN1(n5613),
    .DIN1_t(n5613_t),
    .DIN2(n3866),
    .DIN2_t(n3866_t),
    .Q(n3865),
    .Q_t(n3865_t)
  );


  xor2s3
  U2345
  (
    .DIN1(n5611),
    .DIN1_t(n5611_t),
    .DIN2(n5612),
    .DIN2_t(n5612_t),
    .Q(n3866),
    .Q_t(n3866_t)
  );


  xor2s3
  U2346
  (
    .DIN1(n5614),
    .DIN1_t(n5614_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3864),
    .Q_t(n3864_t)
  );


  nnd2s3
  U2347
  (
    .DIN1(n3867),
    .DIN1_t(n3867_t),
    .DIN2(n6675),
    .DIN2_t(n6675_t),
    .Q(n3862),
    .Q_t(n3862_t)
  );


  nnd2s3
  U2348
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2105),
    .DIN2_t(n2105_t),
    .Q(n3861),
    .Q_t(n3861_t)
  );


  nnd2s3
  U2349
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2056),
    .DIN2_t(n2056_t),
    .Q(n3860),
    .Q_t(n3860_t)
  );


  nnd4s2
  U2350
  (
    .DIN1(n3868),
    .DIN1_t(n3868_t),
    .DIN2(n3869),
    .DIN2_t(n3869_t),
    .DIN3(n3870),
    .DIN3_t(n3870_t),
    .DIN4(n3871),
    .DIN4_t(n3871_t),
    .Q(WX4535),
    .Q_t(WX4535_t)
  );


  nnd2s3
  U2351
  (
    .DIN1(n3600),
    .DIN1_t(n3600_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3871),
    .Q_t(n3871_t)
  );


  xor2s3
  U2352
  (
    .DIN1(n3872),
    .DIN1_t(n3872_t),
    .DIN2(n3873),
    .DIN2_t(n3873_t),
    .Q(n3600),
    .Q_t(n3600_t)
  );


  xor2s3
  U2353
  (
    .DIN1(n5618),
    .DIN1_t(n5618_t),
    .DIN2(n3874),
    .DIN2_t(n3874_t),
    .Q(n3873),
    .Q_t(n3873_t)
  );


  xor2s3
  U2354
  (
    .DIN1(n5616),
    .DIN1_t(n5616_t),
    .DIN2(n5617),
    .DIN2_t(n5617_t),
    .Q(n3874),
    .Q_t(n3874_t)
  );


  xor2s3
  U2355
  (
    .DIN1(n5619),
    .DIN1_t(n5619_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3872),
    .Q_t(n3872_t)
  );


  nnd2s3
  U2356
  (
    .DIN1(n3875),
    .DIN1_t(n3875_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3870),
    .Q_t(n3870_t)
  );


  nnd2s3
  U2357
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2106),
    .DIN2_t(n2106_t),
    .Q(tempn3869),
    .Q_t(tempn3869_t)
  );


  nnd2s3
  U2358
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2055),
    .DIN2_t(n2055_t),
    .Q(n3868),
    .Q_t(n3868_t)
  );


  nnd4s2
  U2359
  (
    .DIN1(n3876),
    .DIN1_t(n3876_t),
    .DIN2(n3877),
    .DIN2_t(n3877_t),
    .DIN3(n3878),
    .DIN3_t(n3878_t),
    .DIN4(n3879),
    .DIN4_t(n3879_t),
    .Q(WX4533),
    .Q_t(WX4533_t)
  );


  nnd2s3
  U2360
  (
    .DIN1(n3608),
    .DIN1_t(n3608_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3879),
    .Q_t(n3879_t)
  );


  xor2s3
  U2361
  (
    .DIN1(n3880),
    .DIN1_t(n3880_t),
    .DIN2(n3881),
    .DIN2_t(n3881_t),
    .Q(n3608),
    .Q_t(n3608_t)
  );


  xor2s3
  U2362
  (
    .DIN1(n5623),
    .DIN1_t(n5623_t),
    .DIN2(n3882),
    .DIN2_t(n3882_t),
    .Q(n3881),
    .Q_t(n3881_t)
  );


  xor2s3
  U2363
  (
    .DIN1(n5621),
    .DIN1_t(n5621_t),
    .DIN2(n5622),
    .DIN2_t(n5622_t),
    .Q(n3882),
    .Q_t(n3882_t)
  );


  xor2s3
  U2364
  (
    .DIN1(n5624),
    .DIN1_t(n5624_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3880),
    .Q_t(n3880_t)
  );


  nnd2s3
  U2365
  (
    .DIN1(n3883),
    .DIN1_t(n3883_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3878),
    .Q_t(n3878_t)
  );


  nnd2s3
  U2366
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2107),
    .DIN2_t(n2107_t),
    .Q(n3877),
    .Q_t(n3877_t)
  );


  nnd2s3
  U2367
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2054),
    .DIN2_t(n2054_t),
    .Q(n3876),
    .Q_t(n3876_t)
  );


  nnd4s2
  U2368
  (
    .DIN1(n3884),
    .DIN1_t(n3884_t),
    .DIN2(n3885),
    .DIN2_t(n3885_t),
    .DIN3(n3886),
    .DIN3_t(n3886_t),
    .DIN4(n3887),
    .DIN4_t(n3887_t),
    .Q(WX4531),
    .Q_t(WX4531_t)
  );


  nnd2s3
  U2369
  (
    .DIN1(n3616),
    .DIN1_t(n3616_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3887),
    .Q_t(n3887_t)
  );


  xor2s3
  U2370
  (
    .DIN1(n3888),
    .DIN1_t(n3888_t),
    .DIN2(n3889),
    .DIN2_t(n3889_t),
    .Q(n3616),
    .Q_t(n3616_t)
  );


  xor2s3
  U2371
  (
    .DIN1(n5628),
    .DIN1_t(n5628_t),
    .DIN2(n3890),
    .DIN2_t(n3890_t),
    .Q(n3889),
    .Q_t(n3889_t)
  );


  xor2s3
  U2372
  (
    .DIN1(n5626),
    .DIN1_t(n5626_t),
    .DIN2(n5627),
    .DIN2_t(n5627_t),
    .Q(n3890),
    .Q_t(n3890_t)
  );


  xor2s3
  U2373
  (
    .DIN1(n5629),
    .DIN1_t(n5629_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3888),
    .Q_t(n3888_t)
  );


  nnd2s3
  U2374
  (
    .DIN1(n3891),
    .DIN1_t(n3891_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3886),
    .Q_t(n3886_t)
  );


  nnd2s3
  U2375
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2108),
    .DIN2_t(n2108_t),
    .Q(n3885),
    .Q_t(n3885_t)
  );


  nnd2s3
  U2376
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2053),
    .DIN2_t(n2053_t),
    .Q(n3884),
    .Q_t(n3884_t)
  );


  nnd4s2
  U2377
  (
    .DIN1(n3892),
    .DIN1_t(n3892_t),
    .DIN2(n3893),
    .DIN2_t(n3893_t),
    .DIN3(n3894),
    .DIN3_t(n3894_t),
    .DIN4(n3895),
    .DIN4_t(n3895_t),
    .Q(WX4529),
    .Q_t(WX4529_t)
  );


  nnd2s3
  U2378
  (
    .DIN1(n3624),
    .DIN1_t(n3624_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3895),
    .Q_t(n3895_t)
  );


  xor2s3
  U2379
  (
    .DIN1(n3896),
    .DIN1_t(n3896_t),
    .DIN2(n3897),
    .DIN2_t(n3897_t),
    .Q(n3624),
    .Q_t(n3624_t)
  );


  xor2s3
  U2380
  (
    .DIN1(n5633),
    .DIN1_t(n5633_t),
    .DIN2(n3898),
    .DIN2_t(n3898_t),
    .Q(n3897),
    .Q_t(n3897_t)
  );


  xor2s3
  U2381
  (
    .DIN1(n5631),
    .DIN1_t(n5631_t),
    .DIN2(n5632),
    .DIN2_t(n5632_t),
    .Q(n3898),
    .Q_t(n3898_t)
  );


  xor2s3
  U2382
  (
    .DIN1(n5634),
    .DIN1_t(n5634_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3896),
    .Q_t(n3896_t)
  );


  nnd2s3
  U2383
  (
    .DIN1(n3899),
    .DIN1_t(n3899_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3894),
    .Q_t(n3894_t)
  );


  nnd2s3
  U2384
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2109),
    .DIN2_t(n2109_t),
    .Q(n3893),
    .Q_t(n3893_t)
  );


  nnd2s3
  U2385
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2052),
    .DIN2_t(n2052_t),
    .Q(n3892),
    .Q_t(n3892_t)
  );


  nnd4s2
  U2386
  (
    .DIN1(n3900),
    .DIN1_t(n3900_t),
    .DIN2(n3901),
    .DIN2_t(n3901_t),
    .DIN3(n3902),
    .DIN3_t(n3902_t),
    .DIN4(n3903),
    .DIN4_t(n3903_t),
    .Q(WX4527),
    .Q_t(WX4527_t)
  );


  nnd2s3
  U2387
  (
    .DIN1(n3632),
    .DIN1_t(n3632_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3903),
    .Q_t(n3903_t)
  );


  xor2s3
  U2388
  (
    .DIN1(n3904),
    .DIN1_t(n3904_t),
    .DIN2(n3905),
    .DIN2_t(n3905_t),
    .Q(n3632),
    .Q_t(n3632_t)
  );


  xor2s3
  U2389
  (
    .DIN1(n5638),
    .DIN1_t(n5638_t),
    .DIN2(n3906),
    .DIN2_t(n3906_t),
    .Q(n3905),
    .Q_t(n3905_t)
  );


  xor2s3
  U2390
  (
    .DIN1(n5636),
    .DIN1_t(n5636_t),
    .DIN2(n5637),
    .DIN2_t(n5637_t),
    .Q(n3906),
    .Q_t(n3906_t)
  );


  xor2s3
  U2391
  (
    .DIN1(n5639),
    .DIN1_t(n5639_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3904),
    .Q_t(n3904_t)
  );


  nnd2s3
  U2392
  (
    .DIN1(n3907),
    .DIN1_t(n3907_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3902),
    .Q_t(n3902_t)
  );


  nnd2s3
  U2393
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2110),
    .DIN2_t(n2110_t),
    .Q(n3901),
    .Q_t(n3901_t)
  );


  nnd2s3
  U2394
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2051),
    .DIN2_t(n2051_t),
    .Q(n3900),
    .Q_t(n3900_t)
  );


  nnd4s2
  U2395
  (
    .DIN1(n3908),
    .DIN1_t(n3908_t),
    .DIN2(n3909),
    .DIN2_t(n3909_t),
    .DIN3(n3910),
    .DIN3_t(n3910_t),
    .DIN4(n3911),
    .DIN4_t(n3911_t),
    .Q(WX4525),
    .Q_t(WX4525_t)
  );


  nnd2s3
  U2396
  (
    .DIN1(n3640),
    .DIN1_t(n3640_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3911),
    .Q_t(n3911_t)
  );


  xor2s3
  U2397
  (
    .DIN1(n3912),
    .DIN1_t(n3912_t),
    .DIN2(n3913),
    .DIN2_t(n3913_t),
    .Q(n3640),
    .Q_t(n3640_t)
  );


  xor2s3
  U2398
  (
    .DIN1(n5643),
    .DIN1_t(n5643_t),
    .DIN2(n3914),
    .DIN2_t(n3914_t),
    .Q(n3913),
    .Q_t(n3913_t)
  );


  xor2s3
  U2399
  (
    .DIN1(n5641),
    .DIN1_t(n5641_t),
    .DIN2(n5642),
    .DIN2_t(n5642_t),
    .Q(n3914),
    .Q_t(n3914_t)
  );


  xor2s3
  U2400
  (
    .DIN1(n5644),
    .DIN1_t(n5644_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3912),
    .Q_t(n3912_t)
  );


  nnd2s3
  U2401
  (
    .DIN1(n3915),
    .DIN1_t(n3915_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3910),
    .Q_t(n3910_t)
  );


  nnd2s3
  U2402
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2111),
    .DIN2_t(n2111_t),
    .Q(n3909),
    .Q_t(n3909_t)
  );


  nnd2s3
  U2403
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2050),
    .DIN2_t(n2050_t),
    .Q(n3908),
    .Q_t(n3908_t)
  );


  nnd4s2
  U2404
  (
    .DIN1(n3916),
    .DIN1_t(n3916_t),
    .DIN2(n3917),
    .DIN2_t(n3917_t),
    .DIN3(n3918),
    .DIN3_t(n3918_t),
    .DIN4(n3919),
    .DIN4_t(n3919_t),
    .Q(WX4523),
    .Q_t(WX4523_t)
  );


  nnd2s3
  U2405
  (
    .DIN1(n3648),
    .DIN1_t(n3648_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3919),
    .Q_t(n3919_t)
  );


  xor2s3
  U2406
  (
    .DIN1(n3920),
    .DIN1_t(n3920_t),
    .DIN2(n3921),
    .DIN2_t(n3921_t),
    .Q(n3648),
    .Q_t(n3648_t)
  );


  xor2s3
  U2407
  (
    .DIN1(n5648),
    .DIN1_t(n5648_t),
    .DIN2(n3922),
    .DIN2_t(n3922_t),
    .Q(n3921),
    .Q_t(n3921_t)
  );


  xor2s3
  U2408
  (
    .DIN1(n5646),
    .DIN1_t(n5646_t),
    .DIN2(n5647),
    .DIN2_t(n5647_t),
    .Q(n3922),
    .Q_t(n3922_t)
  );


  xor2s3
  U2409
  (
    .DIN1(n5649),
    .DIN1_t(n5649_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n3920),
    .Q_t(n3920_t)
  );


  nnd2s3
  U2410
  (
    .DIN1(n3923),
    .DIN1_t(n3923_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3918),
    .Q_t(n3918_t)
  );


  nnd2s3
  U2411
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2112),
    .DIN2_t(n2112_t),
    .Q(n3917),
    .Q_t(n3917_t)
  );


  nnd2s3
  U2412
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2049),
    .DIN2_t(n2049_t),
    .Q(n3916),
    .Q_t(n3916_t)
  );


  nor2s3
  U2413
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n2112),
    .DIN2_t(n2112_t),
    .Q(WX4425),
    .Q_t(WX4425_t)
  );


  nor2s3
  U2414
  (
    .DIN1(n5652),
    .DIN1_t(n5652_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4423),
    .Q_t(WX4423_t)
  );


  nor2s3
  U2415
  (
    .DIN1(n5653),
    .DIN1_t(n5653_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4421),
    .Q_t(WX4421_t)
  );


  nor2s3
  U2416
  (
    .DIN1(n5654),
    .DIN1_t(n5654_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4419),
    .Q_t(WX4419_t)
  );


  nor2s3
  U2417
  (
    .DIN1(n5655),
    .DIN1_t(n5655_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4417),
    .Q_t(WX4417_t)
  );


  nor2s3
  U2418
  (
    .DIN1(n5656),
    .DIN1_t(n5656_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4415),
    .Q_t(WX4415_t)
  );


  nor2s3
  U2419
  (
    .DIN1(n5657),
    .DIN1_t(n5657_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4413),
    .Q_t(WX4413_t)
  );


  nor2s3
  U2420
  (
    .DIN1(n5658),
    .DIN1_t(n5658_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4411),
    .Q_t(WX4411_t)
  );


  nor2s3
  U2421
  (
    .DIN1(n5659),
    .DIN1_t(n5659_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX4409),
    .Q_t(WX4409_t)
  );


  nor2s3
  U2422
  (
    .DIN1(n5660),
    .DIN1_t(n5660_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX4407),
    .Q_t(WX4407_t)
  );


  nor2s3
  U2423
  (
    .DIN1(n5661),
    .DIN1_t(n5661_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX4405),
    .Q_t(WX4405_t)
  );


  nor2s3
  U2424
  (
    .DIN1(n5662),
    .DIN1_t(n5662_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX4403),
    .Q_t(WX4403_t)
  );


  nor2s3
  U2425
  (
    .DIN1(n5663),
    .DIN1_t(n5663_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX4401),
    .Q_t(WX4401_t)
  );


  nor2s3
  U2426
  (
    .DIN1(n5664),
    .DIN1_t(n5664_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX4399),
    .Q_t(WX4399_t)
  );


  nor2s3
  U2427
  (
    .DIN1(n5665),
    .DIN1_t(n5665_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX4397),
    .Q_t(WX4397_t)
  );


  nor2s3
  U2428
  (
    .DIN1(n5666),
    .DIN1_t(n5666_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX4395),
    .Q_t(WX4395_t)
  );


  nor2s3
  U2429
  (
    .DIN1(n5667),
    .DIN1_t(n5667_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX4393),
    .Q_t(WX4393_t)
  );


  nor2s3
  U2430
  (
    .DIN1(n5668),
    .DIN1_t(n5668_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX4391),
    .Q_t(WX4391_t)
  );


  nor2s3
  U2431
  (
    .DIN1(n5669),
    .DIN1_t(n5669_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX4389),
    .Q_t(WX4389_t)
  );


  nor2s3
  U2432
  (
    .DIN1(n5670),
    .DIN1_t(n5670_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX4387),
    .Q_t(WX4387_t)
  );


  nor2s3
  U2433
  (
    .DIN1(n5671),
    .DIN1_t(n5671_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4385),
    .Q_t(WX4385_t)
  );


  nor2s3
  U2434
  (
    .DIN1(n5672),
    .DIN1_t(n5672_t),
    .DIN2(n6777),
    .DIN2_t(n6777_t),
    .Q(WX4383),
    .Q_t(WX4383_t)
  );


  nor2s3
  U2435
  (
    .DIN1(n5673),
    .DIN1_t(n5673_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4381),
    .Q_t(WX4381_t)
  );


  nor2s3
  U2436
  (
    .DIN1(n5674),
    .DIN1_t(n5674_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4379),
    .Q_t(WX4379_t)
  );


  nor2s3
  U2437
  (
    .DIN1(n5675),
    .DIN1_t(n5675_t),
    .DIN2(n6778),
    .DIN2_t(n6778_t),
    .Q(WX4377),
    .Q_t(WX4377_t)
  );


  nor2s3
  U2438
  (
    .DIN1(n5676),
    .DIN1_t(n5676_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX4375),
    .Q_t(WX4375_t)
  );


  nor2s3
  U2439
  (
    .DIN1(n5677),
    .DIN1_t(n5677_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX4373),
    .Q_t(WX4373_t)
  );


  nor2s3
  U2440
  (
    .DIN1(n5678),
    .DIN1_t(n5678_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX4371),
    .Q_t(WX4371_t)
  );


  nor2s3
  U2441
  (
    .DIN1(n5679),
    .DIN1_t(n5679_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX4369),
    .Q_t(WX4369_t)
  );


  nor2s3
  U2442
  (
    .DIN1(n5680),
    .DIN1_t(n5680_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX4367),
    .Q_t(WX4367_t)
  );


  nor2s3
  U2443
  (
    .DIN1(n5681),
    .DIN1_t(n5681_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX4365),
    .Q_t(WX4365_t)
  );


  nor2s3
  U2444
  (
    .DIN1(n5682),
    .DIN1_t(n5682_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX4363),
    .Q_t(WX4363_t)
  );


  nor2s3
  U2445
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3924),
    .DIN2_t(n3924_t),
    .Q(WX3912),
    .Q_t(WX3912_t)
  );


  xor2s3
  U2446
  (
    .DIN1(n5821),
    .DIN1_t(n5821_t),
    .DIN2(n6109),
    .DIN2_t(n6109_t),
    .Q(n3924),
    .Q_t(n3924_t)
  );


  nor2s3
  U2447
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3925),
    .DIN2_t(n3925_t),
    .Q(WX3910),
    .Q_t(WX3910_t)
  );


  xor2s3
  U2448
  (
    .DIN1(n5816),
    .DIN1_t(n5816_t),
    .DIN2(n6100),
    .DIN2_t(n6100_t),
    .Q(n3925),
    .Q_t(n3925_t)
  );


  nor2s3
  U2449
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3926),
    .DIN2_t(n3926_t),
    .Q(WX3908),
    .Q_t(WX3908_t)
  );


  xor2s3
  U2450
  (
    .DIN1(n5811),
    .DIN1_t(n5811_t),
    .DIN2(n6091),
    .DIN2_t(n6091_t),
    .Q(n3926),
    .Q_t(n3926_t)
  );


  nor2s3
  U2451
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3927),
    .DIN2_t(n3927_t),
    .Q(WX3906),
    .Q_t(WX3906_t)
  );


  xor2s3
  U2452
  (
    .DIN1(n5806),
    .DIN1_t(n5806_t),
    .DIN2(n6082),
    .DIN2_t(n6082_t),
    .Q(n3927),
    .Q_t(n3927_t)
  );


  nor2s3
  U2453
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3928),
    .DIN2_t(n3928_t),
    .Q(WX3904),
    .Q_t(WX3904_t)
  );


  xor2s3
  U2454
  (
    .DIN1(n5801),
    .DIN1_t(n5801_t),
    .DIN2(n6073),
    .DIN2_t(n6073_t),
    .Q(n3928),
    .Q_t(n3928_t)
  );


  nor2s3
  U2455
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3929),
    .DIN2_t(n3929_t),
    .Q(WX3902),
    .Q_t(WX3902_t)
  );


  xor2s3
  U2456
  (
    .DIN1(n5796),
    .DIN1_t(n5796_t),
    .DIN2(n6064),
    .DIN2_t(n6064_t),
    .Q(n3929),
    .Q_t(n3929_t)
  );


  nor2s3
  U2457
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3930),
    .DIN2_t(n3930_t),
    .Q(WX3900),
    .Q_t(WX3900_t)
  );


  xor2s3
  U2458
  (
    .DIN1(n5791),
    .DIN1_t(n5791_t),
    .DIN2(n6055),
    .DIN2_t(n6055_t),
    .Q(n3930),
    .Q_t(n3930_t)
  );


  nor2s3
  U2459
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3931),
    .DIN2_t(n3931_t),
    .Q(WX3898),
    .Q_t(WX3898_t)
  );


  xor2s3
  U2460
  (
    .DIN1(n5786),
    .DIN1_t(n5786_t),
    .DIN2(n6046),
    .DIN2_t(n6046_t),
    .Q(n3931),
    .Q_t(n3931_t)
  );


  nor2s3
  U2461
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3932),
    .DIN2_t(n3932_t),
    .Q(WX3896),
    .Q_t(WX3896_t)
  );


  xor2s3
  U2462
  (
    .DIN1(n5781),
    .DIN1_t(n5781_t),
    .DIN2(n6037),
    .DIN2_t(n6037_t),
    .Q(n3932),
    .Q_t(n3932_t)
  );


  nor2s3
  U2463
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3933),
    .DIN2_t(n3933_t),
    .Q(WX3894),
    .Q_t(WX3894_t)
  );


  xor2s3
  U2464
  (
    .DIN1(n5776),
    .DIN1_t(n5776_t),
    .DIN2(n6028),
    .DIN2_t(n6028_t),
    .Q(n3933),
    .Q_t(n3933_t)
  );


  nor2s3
  U2465
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3934),
    .DIN2_t(n3934_t),
    .Q(WX3892),
    .Q_t(WX3892_t)
  );


  xor2s3
  U2466
  (
    .DIN1(n5771),
    .DIN1_t(n5771_t),
    .DIN2(n6019),
    .DIN2_t(n6019_t),
    .Q(n3934),
    .Q_t(n3934_t)
  );


  nor2s3
  U2467
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3935),
    .DIN2_t(n3935_t),
    .Q(WX3890),
    .Q_t(WX3890_t)
  );


  xor2s3
  U2468
  (
    .DIN1(n5766),
    .DIN1_t(n5766_t),
    .DIN2(n6010),
    .DIN2_t(n6010_t),
    .Q(n3935),
    .Q_t(n3935_t)
  );


  nor2s3
  U2469
  (
    .DIN1(n6804),
    .DIN1_t(n6804_t),
    .DIN2(n3936),
    .DIN2_t(n3936_t),
    .Q(WX3888),
    .Q_t(WX3888_t)
  );


  xor2s3
  U2470
  (
    .DIN1(n5761),
    .DIN1_t(n5761_t),
    .DIN2(n6001),
    .DIN2_t(n6001_t),
    .Q(n3936),
    .Q_t(n3936_t)
  );


  nor2s3
  U2471
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3937),
    .DIN2_t(n3937_t),
    .Q(WX3886),
    .Q_t(WX3886_t)
  );


  xor2s3
  U2472
  (
    .DIN1(n5756),
    .DIN1_t(n5756_t),
    .DIN2(n5992),
    .DIN2_t(n5992_t),
    .Q(n3937),
    .Q_t(n3937_t)
  );


  nor2s3
  U2473
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3938),
    .DIN2_t(n3938_t),
    .Q(WX3884),
    .Q_t(WX3884_t)
  );


  xor2s3
  U2474
  (
    .DIN1(n5751),
    .DIN1_t(n5751_t),
    .DIN2(n5983),
    .DIN2_t(n5983_t),
    .Q(n3938),
    .Q_t(n3938_t)
  );


  nor2s3
  U2475
  (
    .DIN1(n3939),
    .DIN1_t(n3939_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX3882),
    .Q_t(WX3882_t)
  );


  xnr2s3
  U2476
  (
    .DIN1(n5974),
    .DIN1_t(n5974_t),
    .DIN2(n3940),
    .DIN2_t(n3940_t),
    .Q(n3939),
    .Q_t(n3939_t)
  );


  xor2s3
  U2477
  (
    .DIN1(n5746),
    .DIN1_t(n5746_t),
    .DIN2(n5826),
    .DIN2_t(n5826_t),
    .Q(n3940),
    .Q_t(n3940_t)
  );


  nor2s3
  U2478
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3941),
    .DIN2_t(n3941_t),
    .Q(WX3880),
    .Q_t(WX3880_t)
  );


  xor2s3
  U2479
  (
    .DIN1(n5742),
    .DIN1_t(n5742_t),
    .DIN2(n3315),
    .DIN2_t(n3315_t),
    .Q(n3941),
    .Q_t(n3941_t)
  );


  nor2s3
  U2480
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3942),
    .DIN2_t(n3942_t),
    .Q(WX3878),
    .Q_t(WX3878_t)
  );


  xor2s3
  U2481
  (
    .DIN1(n5738),
    .DIN1_t(n5738_t),
    .DIN2(n3313),
    .DIN2_t(n3313_t),
    .Q(n3942),
    .Q_t(n3942_t)
  );


  nor2s3
  U2482
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3943),
    .DIN2_t(n3943_t),
    .Q(WX3876),
    .Q_t(WX3876_t)
  );


  xor2s3
  U2483
  (
    .DIN1(n5734),
    .DIN1_t(n5734_t),
    .DIN2(n3311),
    .DIN2_t(n3311_t),
    .Q(n3943),
    .Q_t(n3943_t)
  );


  nor2s3
  U2484
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3944),
    .DIN2_t(n3944_t),
    .Q(WX3874),
    .Q_t(WX3874_t)
  );


  xor2s3
  U2485
  (
    .DIN1(n5730),
    .DIN1_t(n5730_t),
    .DIN2(n3309),
    .DIN2_t(n3309_t),
    .Q(n3944),
    .Q_t(n3944_t)
  );


  nor2s3
  U2486
  (
    .DIN1(n3945),
    .DIN1_t(n3945_t),
    .DIN2(n6779),
    .DIN2_t(n6779_t),
    .Q(WX3872),
    .Q_t(WX3872_t)
  );


  xnr2s3
  U2487
  (
    .DIN1(n3307),
    .DIN1_t(n3307_t),
    .DIN2(n3946),
    .DIN2_t(n3946_t),
    .Q(n3945),
    .Q_t(n3945_t)
  );


  xor2s3
  U2488
  (
    .DIN1(n5726),
    .DIN1_t(n5726_t),
    .DIN2(n5826),
    .DIN2_t(n5826_t),
    .Q(n3946),
    .Q_t(n3946_t)
  );


  nor2s3
  U2489
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3947),
    .DIN2_t(n3947_t),
    .Q(WX3870),
    .Q_t(WX3870_t)
  );


  xor2s3
  U2490
  (
    .DIN1(n5722),
    .DIN1_t(n5722_t),
    .DIN2(n3305),
    .DIN2_t(n3305_t),
    .Q(n3947),
    .Q_t(n3947_t)
  );


  nor2s3
  U2491
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3948),
    .DIN2_t(n3948_t),
    .Q(WX3868),
    .Q_t(WX3868_t)
  );


  xor2s3
  U2492
  (
    .DIN1(n5718),
    .DIN1_t(n5718_t),
    .DIN2(n3303),
    .DIN2_t(n3303_t),
    .Q(n3948),
    .Q_t(n3948_t)
  );


  nor2s3
  U2493
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3949),
    .DIN2_t(n3949_t),
    .Q(WX3866),
    .Q_t(WX3866_t)
  );


  xor2s3
  U2494
  (
    .DIN1(n5714),
    .DIN1_t(n5714_t),
    .DIN2(n3301),
    .DIN2_t(n3301_t),
    .Q(n3949),
    .Q_t(n3949_t)
  );


  nor2s3
  U2495
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3950),
    .DIN2_t(n3950_t),
    .Q(WX3864),
    .Q_t(WX3864_t)
  );


  xor2s3
  U2496
  (
    .DIN1(n5710),
    .DIN1_t(n5710_t),
    .DIN2(n3299),
    .DIN2_t(n3299_t),
    .Q(n3950),
    .Q_t(n3950_t)
  );


  nor2s3
  U2497
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3951),
    .DIN2_t(n3951_t),
    .Q(WX3862),
    .Q_t(WX3862_t)
  );


  xor2s3
  U2498
  (
    .DIN1(n5706),
    .DIN1_t(n5706_t),
    .DIN2(n3297),
    .DIN2_t(n3297_t),
    .Q(n3951),
    .Q_t(n3951_t)
  );


  nor2s3
  U2499
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n3952),
    .DIN2_t(n3952_t),
    .Q(WX3860),
    .Q_t(WX3860_t)
  );


  xor2s3
  U2500
  (
    .DIN1(n5702),
    .DIN1_t(n5702_t),
    .DIN2(n3295),
    .DIN2_t(n3295_t),
    .Q(n3952),
    .Q_t(n3952_t)
  );


  nor2s3
  U2501
  (
    .DIN1(n3953),
    .DIN1_t(n3953_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX3858),
    .Q_t(WX3858_t)
  );


  xnr2s3
  U2502
  (
    .DIN1(n3293),
    .DIN1_t(n3293_t),
    .DIN2(n3954),
    .DIN2_t(n3954_t),
    .Q(n3953),
    .Q_t(n3953_t)
  );


  xor2s3
  U2503
  (
    .DIN1(n5698),
    .DIN1_t(n5698_t),
    .DIN2(n5826),
    .DIN2_t(n5826_t),
    .Q(n3954),
    .Q_t(n3954_t)
  );


  nor2s3
  U2504
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n3955),
    .DIN2_t(n3955_t),
    .Q(WX3856),
    .Q_t(WX3856_t)
  );


  xor2s3
  U2505
  (
    .DIN1(n5694),
    .DIN1_t(n5694_t),
    .DIN2(n3291),
    .DIN2_t(n3291_t),
    .Q(n3955),
    .Q_t(n3955_t)
  );


  nor2s3
  U2506
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n3956),
    .DIN2_t(n3956_t),
    .Q(WX3854),
    .Q_t(WX3854_t)
  );


  xor2s3
  U2507
  (
    .DIN1(n5690),
    .DIN1_t(n5690_t),
    .DIN2(n3289),
    .DIN2_t(n3289_t),
    .Q(n3956),
    .Q_t(n3956_t)
  );


  nor2s3
  U2508
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n3957),
    .DIN2_t(n3957_t),
    .Q(WX3852),
    .Q_t(WX3852_t)
  );


  xor2s3
  U2509
  (
    .DIN1(n5686),
    .DIN1_t(n5686_t),
    .DIN2(n3287),
    .DIN2_t(n3287_t),
    .Q(n3957),
    .Q_t(n3957_t)
  );


  nor2s3
  U2510
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n3958),
    .DIN2_t(n3958_t),
    .Q(WX3850),
    .Q_t(WX3850_t)
  );


  xor2s3
  U2511
  (
    .DIN1(n5826),
    .DIN1_t(n5826_t),
    .DIN2(n3285),
    .DIN2_t(n3285_t),
    .Q(n3958),
    .Q_t(n3958_t)
  );


  nor2s3
  U2512
  (
    .DIN1(n5861),
    .DIN1_t(n5861_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX3484),
    .Q_t(WX3484_t)
  );


  nor2s3
  U2513
  (
    .DIN1(n5868),
    .DIN1_t(n5868_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX3482),
    .Q_t(WX3482_t)
  );


  nor2s3
  U2514
  (
    .DIN1(n5875),
    .DIN1_t(n5875_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX3480),
    .Q_t(WX3480_t)
  );


  nor2s3
  U2515
  (
    .DIN1(n5882),
    .DIN1_t(n5882_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX3478),
    .Q_t(WX3478_t)
  );


  nor2s3
  U2516
  (
    .DIN1(n5889),
    .DIN1_t(n5889_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX3476),
    .Q_t(WX3476_t)
  );


  nor2s3
  U2517
  (
    .DIN1(n5896),
    .DIN1_t(n5896_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX3474),
    .Q_t(WX3474_t)
  );


  nor2s3
  U2518
  (
    .DIN1(n5903),
    .DIN1_t(n5903_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX3472),
    .Q_t(WX3472_t)
  );


  nor2s3
  U2519
  (
    .DIN1(n5910),
    .DIN1_t(n5910_t),
    .DIN2(n6780),
    .DIN2_t(n6780_t),
    .Q(WX3470),
    .Q_t(WX3470_t)
  );


  nor2s3
  U2520
  (
    .DIN1(n5917),
    .DIN1_t(n5917_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX3468),
    .Q_t(WX3468_t)
  );


  nor2s3
  U2521
  (
    .DIN1(n5924),
    .DIN1_t(n5924_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX3466),
    .Q_t(WX3466_t)
  );


  nor2s3
  U2522
  (
    .DIN1(n5931),
    .DIN1_t(n5931_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX3464),
    .Q_t(WX3464_t)
  );


  nor2s3
  U2523
  (
    .DIN1(n5938),
    .DIN1_t(n5938_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX3462),
    .Q_t(WX3462_t)
  );


  nor2s3
  U2524
  (
    .DIN1(n5945),
    .DIN1_t(n5945_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX3460),
    .Q_t(WX3460_t)
  );


  nor2s3
  U2525
  (
    .DIN1(n5952),
    .DIN1_t(n5952_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX3458),
    .Q_t(WX3458_t)
  );


  nor2s3
  U2526
  (
    .DIN1(n5959),
    .DIN1_t(n5959_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX3456),
    .Q_t(WX3456_t)
  );


  nor2s3
  U2527
  (
    .DIN1(n5966),
    .DIN1_t(n5966_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX3454),
    .Q_t(WX3454_t)
  );


  nor2s3
  U2528
  (
    .DIN1(n5973),
    .DIN1_t(n5973_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX3452),
    .Q_t(WX3452_t)
  );


  nor2s3
  U2529
  (
    .DIN1(n5982),
    .DIN1_t(n5982_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX3450),
    .Q_t(WX3450_t)
  );


  nor2s3
  U2530
  (
    .DIN1(n5991),
    .DIN1_t(n5991_t),
    .DIN2(n6781),
    .DIN2_t(n6781_t),
    .Q(WX3448),
    .Q_t(WX3448_t)
  );


  nor2s3
  U2531
  (
    .DIN1(n6000),
    .DIN1_t(n6000_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX3446),
    .Q_t(WX3446_t)
  );


  nor2s3
  U2532
  (
    .DIN1(n6009),
    .DIN1_t(n6009_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX3444),
    .Q_t(WX3444_t)
  );


  nor2s3
  U2533
  (
    .DIN1(n6018),
    .DIN1_t(n6018_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX3442),
    .Q_t(WX3442_t)
  );


  nor2s3
  U2534
  (
    .DIN1(n6027),
    .DIN1_t(n6027_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX3440),
    .Q_t(WX3440_t)
  );


  nor2s3
  U2535
  (
    .DIN1(n6036),
    .DIN1_t(n6036_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX3438),
    .Q_t(WX3438_t)
  );


  nor2s3
  U2536
  (
    .DIN1(n6045),
    .DIN1_t(n6045_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX3436),
    .Q_t(WX3436_t)
  );


  nor2s3
  U2537
  (
    .DIN1(n6054),
    .DIN1_t(n6054_t),
    .DIN2(n6782),
    .DIN2_t(n6782_t),
    .Q(WX3434),
    .Q_t(WX3434_t)
  );


  nor2s3
  U2538
  (
    .DIN1(n6063),
    .DIN1_t(n6063_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX3432),
    .Q_t(WX3432_t)
  );


  nor2s3
  U2539
  (
    .DIN1(n6072),
    .DIN1_t(n6072_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX3430),
    .Q_t(WX3430_t)
  );


  nor2s3
  U2540
  (
    .DIN1(n6081),
    .DIN1_t(n6081_t),
    .DIN2(n6787),
    .DIN2_t(n6787_t),
    .Q(WX3428),
    .Q_t(WX3428_t)
  );


  nor2s3
  U2541
  (
    .DIN1(n6090),
    .DIN1_t(n6090_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX3426),
    .Q_t(WX3426_t)
  );


  nor2s3
  U2542
  (
    .DIN1(n6099),
    .DIN1_t(n6099_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX3424),
    .Q_t(WX3424_t)
  );


  nor2s3
  U2543
  (
    .DIN1(n6108),
    .DIN1_t(n6108_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX3422),
    .Q_t(WX3422_t)
  );


  nor2s3
  U2544
  (
    .DIN1(n5860),
    .DIN1_t(n5860_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX3420),
    .Q_t(WX3420_t)
  );


  nor2s3
  U2545
  (
    .DIN1(n5867),
    .DIN1_t(n5867_t),
    .DIN2(n6786),
    .DIN2_t(n6786_t),
    .Q(WX3418),
    .Q_t(WX3418_t)
  );


  nor2s3
  U2546
  (
    .DIN1(n5874),
    .DIN1_t(n5874_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX3416),
    .Q_t(WX3416_t)
  );


  nor2s3
  U2547
  (
    .DIN1(n5881),
    .DIN1_t(n5881_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX3414),
    .Q_t(WX3414_t)
  );


  nor2s3
  U2548
  (
    .DIN1(n5888),
    .DIN1_t(n5888_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX3412),
    .Q_t(WX3412_t)
  );


  nor2s3
  U2549
  (
    .DIN1(n5895),
    .DIN1_t(n5895_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX3410),
    .Q_t(WX3410_t)
  );


  nor2s3
  U2550
  (
    .DIN1(n5902),
    .DIN1_t(n5902_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX3408),
    .Q_t(WX3408_t)
  );


  nor2s3
  U2551
  (
    .DIN1(n5909),
    .DIN1_t(n5909_t),
    .DIN2(n6785),
    .DIN2_t(n6785_t),
    .Q(WX3406),
    .Q_t(WX3406_t)
  );


  nor2s3
  U2552
  (
    .DIN1(n5916),
    .DIN1_t(n5916_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3404),
    .Q_t(WX3404_t)
  );


  nor2s3
  U2553
  (
    .DIN1(n5923),
    .DIN1_t(n5923_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3402),
    .Q_t(WX3402_t)
  );


  nor2s3
  U2554
  (
    .DIN1(n5930),
    .DIN1_t(n5930_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3400),
    .Q_t(WX3400_t)
  );


  nor2s3
  U2555
  (
    .DIN1(n5937),
    .DIN1_t(n5937_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3398),
    .Q_t(WX3398_t)
  );


  nor2s3
  U2556
  (
    .DIN1(n5944),
    .DIN1_t(n5944_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3396),
    .Q_t(WX3396_t)
  );


  nor2s3
  U2557
  (
    .DIN1(n5951),
    .DIN1_t(n5951_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3394),
    .Q_t(WX3394_t)
  );


  nor2s3
  U2558
  (
    .DIN1(n5958),
    .DIN1_t(n5958_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3392),
    .Q_t(WX3392_t)
  );


  nor2s3
  U2559
  (
    .DIN1(n5965),
    .DIN1_t(n5965_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3390),
    .Q_t(WX3390_t)
  );


  and2s3
  U2560
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5972),
    .DIN2_t(n5972_t),
    .Q(WX3388),
    .Q_t(WX3388_t)
  );


  and2s3
  U2561
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5981),
    .DIN2_t(n5981_t),
    .Q(WX3386),
    .Q_t(WX3386_t)
  );


  and2s3
  U2562
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5990),
    .DIN2_t(n5990_t),
    .Q(WX3384),
    .Q_t(WX3384_t)
  );


  and2s3
  U2563
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5999),
    .DIN2_t(n5999_t),
    .Q(WX3382),
    .Q_t(WX3382_t)
  );


  and2s3
  U2564
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6008),
    .DIN2_t(n6008_t),
    .Q(WX3380),
    .Q_t(WX3380_t)
  );


  and2s3
  U2565
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6017),
    .DIN2_t(n6017_t),
    .Q(WX3378),
    .Q_t(WX3378_t)
  );


  and2s3
  U2566
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6026),
    .DIN2_t(n6026_t),
    .Q(WX3376),
    .Q_t(WX3376_t)
  );


  and2s3
  U2567
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6035),
    .DIN2_t(n6035_t),
    .Q(WX3374),
    .Q_t(WX3374_t)
  );


  and2s3
  U2568
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6044),
    .DIN2_t(n6044_t),
    .Q(WX3372),
    .Q_t(WX3372_t)
  );


  and2s3
  U2569
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6053),
    .DIN2_t(n6053_t),
    .Q(WX3370),
    .Q_t(WX3370_t)
  );


  and2s3
  U2570
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6062),
    .DIN2_t(n6062_t),
    .Q(WX3368),
    .Q_t(WX3368_t)
  );


  and2s3
  U2571
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6071),
    .DIN2_t(n6071_t),
    .Q(WX3366),
    .Q_t(WX3366_t)
  );


  and2s3
  U2572
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6080),
    .DIN2_t(n6080_t),
    .Q(WX3364),
    .Q_t(WX3364_t)
  );


  and2s3
  U2573
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6089),
    .DIN2_t(n6089_t),
    .Q(WX3362),
    .Q_t(WX3362_t)
  );


  and2s3
  U2574
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6098),
    .DIN2_t(n6098_t),
    .Q(WX3360),
    .Q_t(WX3360_t)
  );


  and2s3
  U2575
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6107),
    .DIN2_t(n6107_t),
    .Q(WX3358),
    .Q_t(WX3358_t)
  );


  and2s3
  U2576
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5859),
    .DIN2_t(n5859_t),
    .Q(WX3356),
    .Q_t(WX3356_t)
  );


  and2s3
  U2577
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5866),
    .DIN2_t(n5866_t),
    .Q(WX3354),
    .Q_t(WX3354_t)
  );


  and2s3
  U2578
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5873),
    .DIN2_t(n5873_t),
    .Q(WX3352),
    .Q_t(WX3352_t)
  );


  and2s3
  U2579
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5880),
    .DIN2_t(n5880_t),
    .Q(WX3350),
    .Q_t(WX3350_t)
  );


  and2s3
  U2580
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5887),
    .DIN2_t(n5887_t),
    .Q(WX3348),
    .Q_t(WX3348_t)
  );


  and2s3
  U2581
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5894),
    .DIN2_t(n5894_t),
    .Q(WX3346),
    .Q_t(WX3346_t)
  );


  and2s3
  U2582
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5901),
    .DIN2_t(n5901_t),
    .Q(WX3344),
    .Q_t(WX3344_t)
  );


  and2s3
  U2583
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5908),
    .DIN2_t(n5908_t),
    .Q(WX3342),
    .Q_t(WX3342_t)
  );


  and2s3
  U2584
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5915),
    .DIN2_t(n5915_t),
    .Q(WX3340),
    .Q_t(WX3340_t)
  );


  and2s3
  U2585
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5922),
    .DIN2_t(n5922_t),
    .Q(WX3338),
    .Q_t(WX3338_t)
  );


  and2s3
  U2586
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5929),
    .DIN2_t(n5929_t),
    .Q(WX3336),
    .Q_t(WX3336_t)
  );


  and2s3
  U2587
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5936),
    .DIN2_t(n5936_t),
    .Q(WX3334),
    .Q_t(WX3334_t)
  );


  and2s3
  U2588
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5943),
    .DIN2_t(n5943_t),
    .Q(WX3332),
    .Q_t(WX3332_t)
  );


  and2s3
  U2589
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5950),
    .DIN2_t(n5950_t),
    .Q(WX3330),
    .Q_t(WX3330_t)
  );


  and2s3
  U2590
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5957),
    .DIN2_t(n5957_t),
    .Q(WX3328),
    .Q_t(WX3328_t)
  );


  and2s3
  U2591
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5964),
    .DIN2_t(n5964_t),
    .Q(WX3326),
    .Q_t(WX3326_t)
  );


  nor2s3
  U2592
  (
    .DIN1(n5971),
    .DIN1_t(n5971_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3324),
    .Q_t(WX3324_t)
  );


  nor2s3
  U2593
  (
    .DIN1(n5980),
    .DIN1_t(n5980_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3322),
    .Q_t(WX3322_t)
  );


  nor2s3
  U2594
  (
    .DIN1(n5989),
    .DIN1_t(n5989_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3320),
    .Q_t(WX3320_t)
  );


  nor2s3
  U2595
  (
    .DIN1(n5998),
    .DIN1_t(n5998_t),
    .DIN2(n6784),
    .DIN2_t(n6784_t),
    .Q(WX3318),
    .Q_t(WX3318_t)
  );


  nor2s3
  U2596
  (
    .DIN1(n6007),
    .DIN1_t(n6007_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX3316),
    .Q_t(WX3316_t)
  );


  nor2s3
  U2597
  (
    .DIN1(n6016),
    .DIN1_t(n6016_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX3314),
    .Q_t(WX3314_t)
  );


  nor2s3
  U2598
  (
    .DIN1(n6025),
    .DIN1_t(n6025_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX3312),
    .Q_t(WX3312_t)
  );


  nor2s3
  U2599
  (
    .DIN1(n6034),
    .DIN1_t(n6034_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX3310),
    .Q_t(WX3310_t)
  );


  nor2s3
  U2600
  (
    .DIN1(n6043),
    .DIN1_t(n6043_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX3308),
    .Q_t(WX3308_t)
  );


  nor2s3
  U2601
  (
    .DIN1(n6052),
    .DIN1_t(n6052_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX3306),
    .Q_t(WX3306_t)
  );


  nor2s3
  U2602
  (
    .DIN1(n6061),
    .DIN1_t(n6061_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX3304),
    .Q_t(WX3304_t)
  );


  nor2s3
  U2603
  (
    .DIN1(n6070),
    .DIN1_t(n6070_t),
    .DIN2(n6783),
    .DIN2_t(n6783_t),
    .Q(WX3302),
    .Q_t(WX3302_t)
  );


  nor2s3
  U2604
  (
    .DIN1(n6079),
    .DIN1_t(n6079_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX3300),
    .Q_t(WX3300_t)
  );


  nor2s3
  U2605
  (
    .DIN1(n6088),
    .DIN1_t(n6088_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX3298),
    .Q_t(WX3298_t)
  );


  nor2s3
  U2606
  (
    .DIN1(n6097),
    .DIN1_t(n6097_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3296),
    .Q_t(WX3296_t)
  );


  nor2s3
  U2607
  (
    .DIN1(n6106),
    .DIN1_t(n6106_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3294),
    .Q_t(WX3294_t)
  );


  nnd4s2
  U2608
  (
    .DIN1(n3959),
    .DIN1_t(n3959_t),
    .DIN2(n3960),
    .DIN2_t(n3960_t),
    .DIN3(n3961),
    .DIN3_t(n3961_t),
    .DIN4(n3962),
    .DIN4_t(n3962_t),
    .Q(WX3292),
    .Q_t(WX3292_t)
  );


  nnd2s3
  U2609
  (
    .DIN1(n3690),
    .DIN1_t(n3690_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3962),
    .Q_t(n3962_t)
  );


  xor2s3
  U2610
  (
    .DIN1(n3963),
    .DIN1_t(n3963_t),
    .DIN2(n3964),
    .DIN2_t(n3964_t),
    .Q(n3690),
    .Q_t(n3690_t)
  );


  xor2s3
  U2611
  (
    .DIN1(n5683),
    .DIN1_t(n5683_t),
    .DIN2(n5684),
    .DIN2_t(n5684_t),
    .Q(n3964),
    .Q_t(n3964_t)
  );


  xnr2s3
  U2612
  (
    .DIN1(n3269),
    .DIN1_t(n3269_t),
    .DIN2(n5685),
    .DIN2_t(n5685_t),
    .Q(n3963),
    .Q_t(n3963_t)
  );


  nnd2s3
  U2613
  (
    .DIN1(n3965),
    .DIN1_t(n3965_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3961),
    .Q_t(n3961_t)
  );


  nnd2s3
  U2614
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2145),
    .DIN2_t(n2145_t),
    .Q(n3960),
    .Q_t(n3960_t)
  );


  nnd2s3
  U2615
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2144),
    .DIN2_t(n2144_t),
    .Q(n3959),
    .Q_t(n3959_t)
  );


  nnd4s2
  U2616
  (
    .DIN1(n3966),
    .DIN1_t(n3966_t),
    .DIN2(n3967),
    .DIN2_t(n3967_t),
    .DIN3(n3968),
    .DIN3_t(n3968_t),
    .DIN4(n3969),
    .DIN4_t(n3969_t),
    .Q(WX3290),
    .Q_t(WX3290_t)
  );


  nnd2s3
  U2617
  (
    .DIN1(n3697),
    .DIN1_t(n3697_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3969),
    .Q_t(n3969_t)
  );


  xor2s3
  U2618
  (
    .DIN1(n3970),
    .DIN1_t(n3970_t),
    .DIN2(n3971),
    .DIN2_t(n3971_t),
    .Q(n3697),
    .Q_t(n3697_t)
  );


  xor2s3
  U2619
  (
    .DIN1(n5687),
    .DIN1_t(n5687_t),
    .DIN2(n5688),
    .DIN2_t(n5688_t),
    .Q(n3971),
    .Q_t(n3971_t)
  );


  xnr2s3
  U2620
  (
    .DIN1(n3270),
    .DIN1_t(n3270_t),
    .DIN2(n5689),
    .DIN2_t(n5689_t),
    .Q(n3970),
    .Q_t(n3970_t)
  );


  nnd2s3
  U2621
  (
    .DIN1(n3972),
    .DIN1_t(n3972_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3968),
    .Q_t(n3968_t)
  );


  nnd2s3
  U2622
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2146),
    .DIN2_t(n2146_t),
    .Q(n3967),
    .Q_t(n3967_t)
  );


  nnd2s3
  U2623
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2143),
    .DIN2_t(n2143_t),
    .Q(n3966),
    .Q_t(n3966_t)
  );


  nnd4s2
  U2624
  (
    .DIN1(n3973),
    .DIN1_t(n3973_t),
    .DIN2(n3974),
    .DIN2_t(n3974_t),
    .DIN3(n3975),
    .DIN3_t(n3975_t),
    .DIN4(n3976),
    .DIN4_t(n3976_t),
    .Q(WX3288),
    .Q_t(WX3288_t)
  );


  nnd2s3
  U2625
  (
    .DIN1(n3704),
    .DIN1_t(n3704_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3976),
    .Q_t(n3976_t)
  );


  xor2s3
  U2626
  (
    .DIN1(n3977),
    .DIN1_t(n3977_t),
    .DIN2(n3978),
    .DIN2_t(n3978_t),
    .Q(n3704),
    .Q_t(n3704_t)
  );


  xor2s3
  U2627
  (
    .DIN1(n5691),
    .DIN1_t(n5691_t),
    .DIN2(n5692),
    .DIN2_t(n5692_t),
    .Q(n3978),
    .Q_t(n3978_t)
  );


  xnr2s3
  U2628
  (
    .DIN1(n3271),
    .DIN1_t(n3271_t),
    .DIN2(n5693),
    .DIN2_t(n5693_t),
    .Q(n3977),
    .Q_t(n3977_t)
  );


  nnd2s3
  U2629
  (
    .DIN1(n3979),
    .DIN1_t(n3979_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3975),
    .Q_t(n3975_t)
  );


  nnd2s3
  U2630
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2147),
    .DIN2_t(n2147_t),
    .Q(n3974),
    .Q_t(n3974_t)
  );


  nnd2s3
  U2631
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2142),
    .DIN2_t(n2142_t),
    .Q(n3973),
    .Q_t(n3973_t)
  );


  nnd4s2
  U2632
  (
    .DIN1(n3980),
    .DIN1_t(n3980_t),
    .DIN2(n3981),
    .DIN2_t(n3981_t),
    .DIN3(n3982),
    .DIN3_t(n3982_t),
    .DIN4(n3983),
    .DIN4_t(n3983_t),
    .Q(WX3286),
    .Q_t(WX3286_t)
  );


  nnd2s3
  U2633
  (
    .DIN1(n3711),
    .DIN1_t(n3711_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3983),
    .Q_t(n3983_t)
  );


  xor2s3
  U2634
  (
    .DIN1(n3984),
    .DIN1_t(n3984_t),
    .DIN2(n3985),
    .DIN2_t(n3985_t),
    .Q(n3711),
    .Q_t(n3711_t)
  );


  xor2s3
  U2635
  (
    .DIN1(n5695),
    .DIN1_t(n5695_t),
    .DIN2(n5696),
    .DIN2_t(n5696_t),
    .Q(n3985),
    .Q_t(n3985_t)
  );


  xnr2s3
  U2636
  (
    .DIN1(n3272),
    .DIN1_t(n3272_t),
    .DIN2(n5697),
    .DIN2_t(n5697_t),
    .Q(n3984),
    .Q_t(n3984_t)
  );


  nnd2s3
  U2637
  (
    .DIN1(n3986),
    .DIN1_t(n3986_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3982),
    .Q_t(n3982_t)
  );


  nnd2s3
  U2638
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2148),
    .DIN2_t(n2148_t),
    .Q(n3981),
    .Q_t(n3981_t)
  );


  nnd2s3
  U2639
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2141),
    .DIN2_t(n2141_t),
    .Q(n3980),
    .Q_t(n3980_t)
  );


  nnd4s2
  U2640
  (
    .DIN1(n3987),
    .DIN1_t(n3987_t),
    .DIN2(n3988),
    .DIN2_t(n3988_t),
    .DIN3(n3989),
    .DIN3_t(n3989_t),
    .DIN4(n3990),
    .DIN4_t(n3990_t),
    .Q(WX3284),
    .Q_t(WX3284_t)
  );


  nnd2s3
  U2641
  (
    .DIN1(n3718),
    .DIN1_t(n3718_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3990),
    .Q_t(n3990_t)
  );


  xor2s3
  U2642
  (
    .DIN1(n3991),
    .DIN1_t(n3991_t),
    .DIN2(n3992),
    .DIN2_t(n3992_t),
    .Q(n3718),
    .Q_t(n3718_t)
  );


  xor2s3
  U2643
  (
    .DIN1(n5699),
    .DIN1_t(n5699_t),
    .DIN2(n5700),
    .DIN2_t(n5700_t),
    .Q(n3992),
    .Q_t(n3992_t)
  );


  xnr2s3
  U2644
  (
    .DIN1(n3273),
    .DIN1_t(n3273_t),
    .DIN2(n5701),
    .DIN2_t(n5701_t),
    .Q(n3991),
    .Q_t(n3991_t)
  );


  nnd2s3
  U2645
  (
    .DIN1(n3993),
    .DIN1_t(n3993_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3989),
    .Q_t(n3989_t)
  );


  nnd2s3
  U2646
  (
    .DIN1(n6601),
    .DIN1_t(n6601_t),
    .DIN2(n2149),
    .DIN2_t(n2149_t),
    .Q(n3988),
    .Q_t(n3988_t)
  );


  nnd2s3
  U2647
  (
    .DIN1(n6570),
    .DIN1_t(n6570_t),
    .DIN2(n2140),
    .DIN2_t(n2140_t),
    .Q(n3987),
    .Q_t(n3987_t)
  );


  nnd4s2
  U2648
  (
    .DIN1(n3994),
    .DIN1_t(n3994_t),
    .DIN2(n3995),
    .DIN2_t(n3995_t),
    .DIN3(n3996),
    .DIN3_t(n3996_t),
    .DIN4(n3997),
    .DIN4_t(n3997_t),
    .Q(WX3282),
    .Q_t(WX3282_t)
  );


  nnd2s3
  U2649
  (
    .DIN1(n3725),
    .DIN1_t(n3725_t),
    .DIN2(n6643),
    .DIN2_t(n6643_t),
    .Q(n3997),
    .Q_t(n3997_t)
  );


  xor2s3
  U2650
  (
    .DIN1(n3998),
    .DIN1_t(n3998_t),
    .DIN2(n3999),
    .DIN2_t(n3999_t),
    .Q(n3725),
    .Q_t(n3725_t)
  );


  xor2s3
  U2651
  (
    .DIN1(n5703),
    .DIN1_t(n5703_t),
    .DIN2(n5704),
    .DIN2_t(n5704_t),
    .Q(n3999),
    .Q_t(n3999_t)
  );


  xnr2s3
  U2652
  (
    .DIN1(n3274),
    .DIN1_t(n3274_t),
    .DIN2(n5705),
    .DIN2_t(n5705_t),
    .Q(n3998),
    .Q_t(n3998_t)
  );


  nnd2s3
  U2653
  (
    .DIN1(n4000),
    .DIN1_t(n4000_t),
    .DIN2(n6674),
    .DIN2_t(n6674_t),
    .Q(n3996),
    .Q_t(n3996_t)
  );


  nnd2s3
  U2654
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2150),
    .DIN2_t(n2150_t),
    .Q(n3995),
    .Q_t(n3995_t)
  );


  nnd2s3
  U2655
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2139),
    .DIN2_t(n2139_t),
    .Q(n3994),
    .Q_t(n3994_t)
  );


  nnd4s2
  U2656
  (
    .DIN1(n4001),
    .DIN1_t(n4001_t),
    .DIN2(n4002),
    .DIN2_t(n4002_t),
    .DIN3(n4003),
    .DIN3_t(n4003_t),
    .DIN4(n4004),
    .DIN4_t(n4004_t),
    .Q(WX3280),
    .Q_t(WX3280_t)
  );


  nnd2s3
  U2657
  (
    .DIN1(n3732),
    .DIN1_t(n3732_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4004),
    .Q_t(n4004_t)
  );


  xor2s3
  U2658
  (
    .DIN1(n4005),
    .DIN1_t(n4005_t),
    .DIN2(n4006),
    .DIN2_t(n4006_t),
    .Q(n3732),
    .Q_t(n3732_t)
  );


  xor2s3
  U2659
  (
    .DIN1(n5707),
    .DIN1_t(n5707_t),
    .DIN2(n5708),
    .DIN2_t(n5708_t),
    .Q(n4006),
    .Q_t(n4006_t)
  );


  xnr2s3
  U2660
  (
    .DIN1(n3275),
    .DIN1_t(n3275_t),
    .DIN2(n5709),
    .DIN2_t(n5709_t),
    .Q(n4005),
    .Q_t(n4005_t)
  );


  nnd2s3
  U2661
  (
    .DIN1(n4007),
    .DIN1_t(n4007_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4003),
    .Q_t(n4003_t)
  );


  nnd2s3
  U2662
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2151),
    .DIN2_t(n2151_t),
    .Q(n4002),
    .Q_t(n4002_t)
  );


  nnd2s3
  U2663
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2138),
    .DIN2_t(n2138_t),
    .Q(n4001),
    .Q_t(n4001_t)
  );


  nnd4s2
  U2664
  (
    .DIN1(n4008),
    .DIN1_t(n4008_t),
    .DIN2(n4009),
    .DIN2_t(n4009_t),
    .DIN3(n4010),
    .DIN3_t(n4010_t),
    .DIN4(n4011),
    .DIN4_t(n4011_t),
    .Q(WX3278),
    .Q_t(WX3278_t)
  );


  nnd2s3
  U2665
  (
    .DIN1(n3739),
    .DIN1_t(n3739_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4011),
    .Q_t(n4011_t)
  );


  xor2s3
  U2666
  (
    .DIN1(n4012),
    .DIN1_t(n4012_t),
    .DIN2(n4013),
    .DIN2_t(n4013_t),
    .Q(n3739),
    .Q_t(n3739_t)
  );


  xor2s3
  U2667
  (
    .DIN1(n5711),
    .DIN1_t(n5711_t),
    .DIN2(n5712),
    .DIN2_t(n5712_t),
    .Q(n4013),
    .Q_t(n4013_t)
  );


  xnr2s3
  U2668
  (
    .DIN1(n3276),
    .DIN1_t(n3276_t),
    .DIN2(n5713),
    .DIN2_t(n5713_t),
    .Q(n4012),
    .Q_t(n4012_t)
  );


  nnd2s3
  U2669
  (
    .DIN1(n4014),
    .DIN1_t(n4014_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4010),
    .Q_t(n4010_t)
  );


  nnd2s3
  U2670
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2152),
    .DIN2_t(n2152_t),
    .Q(n4009),
    .Q_t(n4009_t)
  );


  nnd2s3
  U2671
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2137),
    .DIN2_t(n2137_t),
    .Q(n4008),
    .Q_t(n4008_t)
  );


  nnd4s2
  U2672
  (
    .DIN1(n4015),
    .DIN1_t(n4015_t),
    .DIN2(n4016),
    .DIN2_t(n4016_t),
    .DIN3(n4017),
    .DIN3_t(n4017_t),
    .DIN4(n4018),
    .DIN4_t(n4018_t),
    .Q(WX3276),
    .Q_t(WX3276_t)
  );


  nnd2s3
  U2673
  (
    .DIN1(n3746),
    .DIN1_t(n3746_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4018),
    .Q_t(n4018_t)
  );


  xor2s3
  U2674
  (
    .DIN1(n4019),
    .DIN1_t(n4019_t),
    .DIN2(n4020),
    .DIN2_t(n4020_t),
    .Q(n3746),
    .Q_t(n3746_t)
  );


  xor2s3
  U2675
  (
    .DIN1(n5715),
    .DIN1_t(n5715_t),
    .DIN2(n5716),
    .DIN2_t(n5716_t),
    .Q(n4020),
    .Q_t(n4020_t)
  );


  xnr2s3
  U2676
  (
    .DIN1(n3277),
    .DIN1_t(n3277_t),
    .DIN2(n5717),
    .DIN2_t(n5717_t),
    .Q(n4019),
    .Q_t(n4019_t)
  );


  nnd2s3
  U2677
  (
    .DIN1(n4021),
    .DIN1_t(n4021_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4017),
    .Q_t(n4017_t)
  );


  nnd2s3
  U2678
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2153),
    .DIN2_t(n2153_t),
    .Q(n4016),
    .Q_t(n4016_t)
  );


  nnd2s3
  U2679
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2136),
    .DIN2_t(n2136_t),
    .Q(n4015),
    .Q_t(n4015_t)
  );


  nnd4s2
  U2680
  (
    .DIN1(n4022),
    .DIN1_t(n4022_t),
    .DIN2(n4023),
    .DIN2_t(n4023_t),
    .DIN3(n4024),
    .DIN3_t(n4024_t),
    .DIN4(n4025),
    .DIN4_t(n4025_t),
    .Q(WX3274),
    .Q_t(WX3274_t)
  );


  nnd2s3
  U2681
  (
    .DIN1(n3753),
    .DIN1_t(n3753_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4025),
    .Q_t(n4025_t)
  );


  xor2s3
  U2682
  (
    .DIN1(n4026),
    .DIN1_t(n4026_t),
    .DIN2(n4027),
    .DIN2_t(n4027_t),
    .Q(n3753),
    .Q_t(n3753_t)
  );


  xor2s3
  U2683
  (
    .DIN1(n5719),
    .DIN1_t(n5719_t),
    .DIN2(n5720),
    .DIN2_t(n5720_t),
    .Q(n4027),
    .Q_t(n4027_t)
  );


  xnr2s3
  U2684
  (
    .DIN1(n3278),
    .DIN1_t(n3278_t),
    .DIN2(n5721),
    .DIN2_t(n5721_t),
    .Q(n4026),
    .Q_t(n4026_t)
  );


  nnd2s3
  U2685
  (
    .DIN1(n4028),
    .DIN1_t(n4028_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4024),
    .Q_t(n4024_t)
  );


  nnd2s3
  U2686
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2154),
    .DIN2_t(n2154_t),
    .Q(n4023),
    .Q_t(n4023_t)
  );


  nnd2s3
  U2687
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2135),
    .DIN2_t(n2135_t),
    .Q(n4022),
    .Q_t(n4022_t)
  );


  nnd4s2
  U2688
  (
    .DIN1(n4029),
    .DIN1_t(n4029_t),
    .DIN2(n4030),
    .DIN2_t(n4030_t),
    .DIN3(n4031),
    .DIN3_t(n4031_t),
    .DIN4(n4032),
    .DIN4_t(n4032_t),
    .Q(WX3272),
    .Q_t(WX3272_t)
  );


  nnd2s3
  U2689
  (
    .DIN1(n3760),
    .DIN1_t(n3760_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4032),
    .Q_t(n4032_t)
  );


  xor2s3
  U2690
  (
    .DIN1(n4033),
    .DIN1_t(n4033_t),
    .DIN2(n4034),
    .DIN2_t(n4034_t),
    .Q(n3760),
    .Q_t(n3760_t)
  );


  xor2s3
  U2691
  (
    .DIN1(n5723),
    .DIN1_t(n5723_t),
    .DIN2(n5724),
    .DIN2_t(n5724_t),
    .Q(n4034),
    .Q_t(n4034_t)
  );


  xnr2s3
  U2692
  (
    .DIN1(n3279),
    .DIN1_t(n3279_t),
    .DIN2(n5725),
    .DIN2_t(n5725_t),
    .Q(n4033),
    .Q_t(n4033_t)
  );


  nnd2s3
  U2693
  (
    .DIN1(n4035),
    .DIN1_t(n4035_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4031),
    .Q_t(n4031_t)
  );


  nnd2s3
  U2694
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2155),
    .DIN2_t(n2155_t),
    .Q(n4030),
    .Q_t(n4030_t)
  );


  nnd2s3
  U2695
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2134),
    .DIN2_t(n2134_t),
    .Q(n4029),
    .Q_t(n4029_t)
  );


  nnd4s2
  U2696
  (
    .DIN1(n4036),
    .DIN1_t(n4036_t),
    .DIN2(n4037),
    .DIN2_t(n4037_t),
    .DIN3(n4038),
    .DIN3_t(n4038_t),
    .DIN4(n4039),
    .DIN4_t(n4039_t),
    .Q(WX3270),
    .Q_t(WX3270_t)
  );


  nnd2s3
  U2697
  (
    .DIN1(n3767),
    .DIN1_t(n3767_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4039),
    .Q_t(n4039_t)
  );


  xor2s3
  U2698
  (
    .DIN1(n4040),
    .DIN1_t(n4040_t),
    .DIN2(n4041),
    .DIN2_t(n4041_t),
    .Q(n3767),
    .Q_t(n3767_t)
  );


  xor2s3
  U2699
  (
    .DIN1(n5727),
    .DIN1_t(n5727_t),
    .DIN2(n5728),
    .DIN2_t(n5728_t),
    .Q(n4041),
    .Q_t(n4041_t)
  );


  xnr2s3
  U2700
  (
    .DIN1(n3280),
    .DIN1_t(n3280_t),
    .DIN2(n5729),
    .DIN2_t(n5729_t),
    .Q(n4040),
    .Q_t(n4040_t)
  );


  nnd2s3
  U2701
  (
    .DIN1(n4042),
    .DIN1_t(n4042_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4038),
    .Q_t(n4038_t)
  );


  nnd2s3
  U2702
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2156),
    .DIN2_t(n2156_t),
    .Q(n4037),
    .Q_t(n4037_t)
  );


  nnd2s3
  U2703
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2133),
    .DIN2_t(n2133_t),
    .Q(n4036),
    .Q_t(n4036_t)
  );


  nnd4s2
  U2704
  (
    .DIN1(n4043),
    .DIN1_t(n4043_t),
    .DIN2(n4044),
    .DIN2_t(n4044_t),
    .DIN3(n4045),
    .DIN3_t(n4045_t),
    .DIN4(n4046),
    .DIN4_t(n4046_t),
    .Q(WX3268),
    .Q_t(WX3268_t)
  );


  nnd2s3
  U2705
  (
    .DIN1(n3774),
    .DIN1_t(n3774_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4046),
    .Q_t(n4046_t)
  );


  xor2s3
  U2706
  (
    .DIN1(n4047),
    .DIN1_t(n4047_t),
    .DIN2(n4048),
    .DIN2_t(n4048_t),
    .Q(n3774),
    .Q_t(n3774_t)
  );


  xor2s3
  U2707
  (
    .DIN1(n5731),
    .DIN1_t(n5731_t),
    .DIN2(n5732),
    .DIN2_t(n5732_t),
    .Q(n4048),
    .Q_t(n4048_t)
  );


  xnr2s3
  U2708
  (
    .DIN1(n3281),
    .DIN1_t(n3281_t),
    .DIN2(n5733),
    .DIN2_t(n5733_t),
    .Q(n4047),
    .Q_t(n4047_t)
  );


  nnd2s3
  U2709
  (
    .DIN1(n4049),
    .DIN1_t(n4049_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4045),
    .Q_t(n4045_t)
  );


  nnd2s3
  U2710
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2157),
    .DIN2_t(n2157_t),
    .Q(n4044),
    .Q_t(n4044_t)
  );


  nnd2s3
  U2711
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2132),
    .DIN2_t(n2132_t),
    .Q(n4043),
    .Q_t(n4043_t)
  );


  nnd4s2
  U2712
  (
    .DIN1(n4050),
    .DIN1_t(n4050_t),
    .DIN2(n4051),
    .DIN2_t(n4051_t),
    .DIN3(n4052),
    .DIN3_t(n4052_t),
    .DIN4(n4053),
    .DIN4_t(n4053_t),
    .Q(WX3266),
    .Q_t(WX3266_t)
  );


  nnd2s3
  U2713
  (
    .DIN1(n3781),
    .DIN1_t(n3781_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4053),
    .Q_t(n4053_t)
  );


  xor2s3
  U2714
  (
    .DIN1(n4054),
    .DIN1_t(n4054_t),
    .DIN2(n4055),
    .DIN2_t(n4055_t),
    .Q(n3781),
    .Q_t(n3781_t)
  );


  xor2s3
  U2715
  (
    .DIN1(n5735),
    .DIN1_t(n5735_t),
    .DIN2(n5736),
    .DIN2_t(n5736_t),
    .Q(n4055),
    .Q_t(n4055_t)
  );


  xnr2s3
  U2716
  (
    .DIN1(n3282),
    .DIN1_t(n3282_t),
    .DIN2(n5737),
    .DIN2_t(n5737_t),
    .Q(n4054),
    .Q_t(n4054_t)
  );


  nnd2s3
  U2717
  (
    .DIN1(n4056),
    .DIN1_t(n4056_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4052),
    .Q_t(n4052_t)
  );


  nnd2s3
  U2718
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2158),
    .DIN2_t(n2158_t),
    .Q(n4051),
    .Q_t(n4051_t)
  );


  nnd2s3
  U2719
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2131),
    .DIN2_t(n2131_t),
    .Q(n4050),
    .Q_t(n4050_t)
  );


  nnd4s2
  U2720
  (
    .DIN1(n4057),
    .DIN1_t(n4057_t),
    .DIN2(n4058),
    .DIN2_t(n4058_t),
    .DIN3(n4059),
    .DIN3_t(n4059_t),
    .DIN4(n4060),
    .DIN4_t(n4060_t),
    .Q(WX3264),
    .Q_t(WX3264_t)
  );


  nnd2s3
  U2721
  (
    .DIN1(n3788),
    .DIN1_t(n3788_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4060),
    .Q_t(n4060_t)
  );


  xor2s3
  U2722
  (
    .DIN1(n4061),
    .DIN1_t(n4061_t),
    .DIN2(n4062),
    .DIN2_t(n4062_t),
    .Q(n3788),
    .Q_t(n3788_t)
  );


  xor2s3
  U2723
  (
    .DIN1(n5739),
    .DIN1_t(n5739_t),
    .DIN2(n5740),
    .DIN2_t(n5740_t),
    .Q(n4062),
    .Q_t(n4062_t)
  );


  xnr2s3
  U2724
  (
    .DIN1(n3283),
    .DIN1_t(n3283_t),
    .DIN2(n5741),
    .DIN2_t(n5741_t),
    .Q(n4061),
    .Q_t(n4061_t)
  );


  nnd2s3
  U2725
  (
    .DIN1(n4063),
    .DIN1_t(n4063_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4059),
    .Q_t(n4059_t)
  );


  nnd2s3
  U2726
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2159),
    .DIN2_t(n2159_t),
    .Q(n4058),
    .Q_t(n4058_t)
  );


  nnd2s3
  U2727
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2130),
    .DIN2_t(n2130_t),
    .Q(n4057),
    .Q_t(n4057_t)
  );


  nnd4s2
  U2728
  (
    .DIN1(n4064),
    .DIN1_t(n4064_t),
    .DIN2(n4065),
    .DIN2_t(n4065_t),
    .DIN3(n4066),
    .DIN3_t(n4066_t),
    .DIN4(n4067),
    .DIN4_t(n4067_t),
    .Q(WX3262),
    .Q_t(WX3262_t)
  );


  nnd2s3
  U2729
  (
    .DIN1(n3795),
    .DIN1_t(n3795_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4067),
    .Q_t(n4067_t)
  );


  xor2s3
  U2730
  (
    .DIN1(n4068),
    .DIN1_t(n4068_t),
    .DIN2(n4069),
    .DIN2_t(n4069_t),
    .Q(n3795),
    .Q_t(n3795_t)
  );


  xor2s3
  U2731
  (
    .DIN1(n5743),
    .DIN1_t(n5743_t),
    .DIN2(n5744),
    .DIN2_t(n5744_t),
    .Q(n4069),
    .Q_t(n4069_t)
  );


  xnr2s3
  U2732
  (
    .DIN1(n3284),
    .DIN1_t(n3284_t),
    .DIN2(n5745),
    .DIN2_t(n5745_t),
    .Q(n4068),
    .Q_t(n4068_t)
  );


  nnd2s3
  U2733
  (
    .DIN1(n4070),
    .DIN1_t(n4070_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4066),
    .Q_t(n4066_t)
  );


  nnd2s3
  U2734
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2160),
    .DIN2_t(n2160_t),
    .Q(n4065),
    .Q_t(n4065_t)
  );


  nnd2s3
  U2735
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2129),
    .DIN2_t(n2129_t),
    .Q(n4064),
    .Q_t(n4064_t)
  );


  nnd4s2
  U2736
  (
    .DIN1(n4071),
    .DIN1_t(n4071_t),
    .DIN2(n4072),
    .DIN2_t(n4072_t),
    .DIN3(n4073),
    .DIN3_t(n4073_t),
    .DIN4(n4074),
    .DIN4_t(n4074_t),
    .Q(WX3260),
    .Q_t(WX3260_t)
  );


  nnd2s3
  U2737
  (
    .DIN1(n3803),
    .DIN1_t(n3803_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4074),
    .Q_t(n4074_t)
  );


  xor2s3
  U2738
  (
    .DIN1(n4075),
    .DIN1_t(n4075_t),
    .DIN2(n4076),
    .DIN2_t(n4076_t),
    .Q(n3803),
    .Q_t(n3803_t)
  );


  xor2s3
  U2739
  (
    .DIN1(n5749),
    .DIN1_t(n5749_t),
    .DIN2(n4077),
    .DIN2_t(n4077_t),
    .Q(n4076),
    .Q_t(n4076_t)
  );


  xor2s3
  U2740
  (
    .DIN1(n5747),
    .DIN1_t(n5747_t),
    .DIN2(n5748),
    .DIN2_t(n5748_t),
    .Q(n4077),
    .Q_t(n4077_t)
  );


  xor2s3
  U2741
  (
    .DIN1(n5750),
    .DIN1_t(n5750_t),
    .DIN2(n6691),
    .DIN2_t(n6691_t),
    .Q(n4075),
    .Q_t(n4075_t)
  );


  nnd2s3
  U2742
  (
    .DIN1(n4078),
    .DIN1_t(n4078_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4073),
    .Q_t(n4073_t)
  );


  nnd2s3
  U2743
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2161),
    .DIN2_t(n2161_t),
    .Q(n4072),
    .Q_t(n4072_t)
  );


  nnd2s3
  U2744
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2128),
    .DIN2_t(n2128_t),
    .Q(n4071),
    .Q_t(n4071_t)
  );


  nnd4s2
  U2745
  (
    .DIN1(n4079),
    .DIN1_t(n4079_t),
    .DIN2(n4080),
    .DIN2_t(n4080_t),
    .DIN3(n4081),
    .DIN3_t(n4081_t),
    .DIN4(n4082),
    .DIN4_t(n4082_t),
    .Q(WX3258),
    .Q_t(WX3258_t)
  );


  nnd2s3
  U2746
  (
    .DIN1(n3811),
    .DIN1_t(n3811_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4082),
    .Q_t(n4082_t)
  );


  xor2s3
  U2747
  (
    .DIN1(n4083),
    .DIN1_t(n4083_t),
    .DIN2(n4084),
    .DIN2_t(n4084_t),
    .Q(n3811),
    .Q_t(n3811_t)
  );


  xor2s3
  U2748
  (
    .DIN1(n5754),
    .DIN1_t(n5754_t),
    .DIN2(n4085),
    .DIN2_t(n4085_t),
    .Q(n4084),
    .Q_t(n4084_t)
  );


  xor2s3
  U2749
  (
    .DIN1(n5752),
    .DIN1_t(n5752_t),
    .DIN2(n5753),
    .DIN2_t(n5753_t),
    .Q(n4085),
    .Q_t(n4085_t)
  );


  xor2s3
  U2750
  (
    .DIN1(n5755),
    .DIN1_t(n5755_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4083),
    .Q_t(n4083_t)
  );


  nnd2s3
  U2751
  (
    .DIN1(n4086),
    .DIN1_t(n4086_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4081),
    .Q_t(n4081_t)
  );


  nnd2s3
  U2752
  (
    .DIN1(n6600),
    .DIN1_t(n6600_t),
    .DIN2(n2162),
    .DIN2_t(n2162_t),
    .Q(n4080),
    .Q_t(n4080_t)
  );


  nnd2s3
  U2753
  (
    .DIN1(n6569),
    .DIN1_t(n6569_t),
    .DIN2(n2127),
    .DIN2_t(n2127_t),
    .Q(n4079),
    .Q_t(n4079_t)
  );


  nnd4s2
  U2754
  (
    .DIN1(n4087),
    .DIN1_t(n4087_t),
    .DIN2(n4088),
    .DIN2_t(n4088_t),
    .DIN3(n4089),
    .DIN3_t(n4089_t),
    .DIN4(n4090),
    .DIN4_t(n4090_t),
    .Q(WX3256),
    .Q_t(WX3256_t)
  );


  nnd2s3
  U2755
  (
    .DIN1(n3819),
    .DIN1_t(n3819_t),
    .DIN2(n6642),
    .DIN2_t(n6642_t),
    .Q(n4090),
    .Q_t(n4090_t)
  );


  xor2s3
  U2756
  (
    .DIN1(n4091),
    .DIN1_t(n4091_t),
    .DIN2(n4092),
    .DIN2_t(n4092_t),
    .Q(n3819),
    .Q_t(n3819_t)
  );


  xor2s3
  U2757
  (
    .DIN1(n5759),
    .DIN1_t(n5759_t),
    .DIN2(n4093),
    .DIN2_t(n4093_t),
    .Q(n4092),
    .Q_t(n4092_t)
  );


  xor2s3
  U2758
  (
    .DIN1(n5757),
    .DIN1_t(n5757_t),
    .DIN2(n5758),
    .DIN2_t(n5758_t),
    .Q(n4093),
    .Q_t(n4093_t)
  );


  xor2s3
  U2759
  (
    .DIN1(n5760),
    .DIN1_t(n5760_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4091),
    .Q_t(n4091_t)
  );


  nnd2s3
  U2760
  (
    .DIN1(n4094),
    .DIN1_t(n4094_t),
    .DIN2(n6673),
    .DIN2_t(n6673_t),
    .Q(n4089),
    .Q_t(n4089_t)
  );


  nnd2s3
  U2761
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2163),
    .DIN2_t(n2163_t),
    .Q(n4088),
    .Q_t(n4088_t)
  );


  nnd2s3
  U2762
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2126),
    .DIN2_t(n2126_t),
    .Q(n4087),
    .Q_t(n4087_t)
  );


  nnd4s2
  U2763
  (
    .DIN1(n4095),
    .DIN1_t(n4095_t),
    .DIN2(n4096),
    .DIN2_t(n4096_t),
    .DIN3(n4097),
    .DIN3_t(n4097_t),
    .DIN4(n4098),
    .DIN4_t(n4098_t),
    .Q(WX3254),
    .Q_t(WX3254_t)
  );


  nnd2s3
  U2764
  (
    .DIN1(n3827),
    .DIN1_t(n3827_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4098),
    .Q_t(n4098_t)
  );


  xor2s3
  U2765
  (
    .DIN1(n4099),
    .DIN1_t(n4099_t),
    .DIN2(n4100),
    .DIN2_t(n4100_t),
    .Q(n3827),
    .Q_t(n3827_t)
  );


  xor2s3
  U2766
  (
    .DIN1(n5764),
    .DIN1_t(n5764_t),
    .DIN2(n4101),
    .DIN2_t(n4101_t),
    .Q(n4100),
    .Q_t(n4100_t)
  );


  xor2s3
  U2767
  (
    .DIN1(n5762),
    .DIN1_t(n5762_t),
    .DIN2(n5763),
    .DIN2_t(n5763_t),
    .Q(n4101),
    .Q_t(n4101_t)
  );


  xor2s3
  U2768
  (
    .DIN1(n5765),
    .DIN1_t(n5765_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4099),
    .Q_t(n4099_t)
  );


  nnd2s3
  U2769
  (
    .DIN1(n4102),
    .DIN1_t(n4102_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4097),
    .Q_t(n4097_t)
  );


  nnd2s3
  U2770
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2164),
    .DIN2_t(n2164_t),
    .Q(n4096),
    .Q_t(n4096_t)
  );


  nnd2s3
  U2771
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2125),
    .DIN2_t(n2125_t),
    .Q(n4095),
    .Q_t(n4095_t)
  );


  nnd4s2
  U2772
  (
    .DIN1(n4103),
    .DIN1_t(n4103_t),
    .DIN2(n4104),
    .DIN2_t(n4104_t),
    .DIN3(n4105),
    .DIN3_t(n4105_t),
    .DIN4(n4106),
    .DIN4_t(n4106_t),
    .Q(WX3252),
    .Q_t(WX3252_t)
  );


  nnd2s3
  U2773
  (
    .DIN1(n3835),
    .DIN1_t(n3835_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4106),
    .Q_t(n4106_t)
  );


  xor2s3
  U2774
  (
    .DIN1(n4107),
    .DIN1_t(n4107_t),
    .DIN2(n4108),
    .DIN2_t(n4108_t),
    .Q(n3835),
    .Q_t(n3835_t)
  );


  xor2s3
  U2775
  (
    .DIN1(n5769),
    .DIN1_t(n5769_t),
    .DIN2(n4109),
    .DIN2_t(n4109_t),
    .Q(n4108),
    .Q_t(n4108_t)
  );


  xor2s3
  U2776
  (
    .DIN1(n5767),
    .DIN1_t(n5767_t),
    .DIN2(n5768),
    .DIN2_t(n5768_t),
    .Q(n4109),
    .Q_t(n4109_t)
  );


  xor2s3
  U2777
  (
    .DIN1(n5770),
    .DIN1_t(n5770_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4107),
    .Q_t(n4107_t)
  );


  nnd2s3
  U2778
  (
    .DIN1(n4110),
    .DIN1_t(n4110_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4105),
    .Q_t(n4105_t)
  );


  nnd2s3
  U2779
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2165),
    .DIN2_t(n2165_t),
    .Q(n4104),
    .Q_t(n4104_t)
  );


  nnd2s3
  U2780
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2124),
    .DIN2_t(n2124_t),
    .Q(n4103),
    .Q_t(n4103_t)
  );


  nnd4s2
  U2781
  (
    .DIN1(n4111),
    .DIN1_t(n4111_t),
    .DIN2(n4112),
    .DIN2_t(n4112_t),
    .DIN3(n4113),
    .DIN3_t(n4113_t),
    .DIN4(n4114),
    .DIN4_t(n4114_t),
    .Q(WX3250),
    .Q_t(WX3250_t)
  );


  nnd2s3
  U2782
  (
    .DIN1(n3843),
    .DIN1_t(n3843_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4114),
    .Q_t(n4114_t)
  );


  xor2s3
  U2783
  (
    .DIN1(n4115),
    .DIN1_t(n4115_t),
    .DIN2(n4116),
    .DIN2_t(n4116_t),
    .Q(n3843),
    .Q_t(n3843_t)
  );


  xor2s3
  U2784
  (
    .DIN1(n5774),
    .DIN1_t(n5774_t),
    .DIN2(n4117),
    .DIN2_t(n4117_t),
    .Q(n4116),
    .Q_t(n4116_t)
  );


  xor2s3
  U2785
  (
    .DIN1(n5772),
    .DIN1_t(n5772_t),
    .DIN2(n5773),
    .DIN2_t(n5773_t),
    .Q(n4117),
    .Q_t(n4117_t)
  );


  xor2s3
  U2786
  (
    .DIN1(n5775),
    .DIN1_t(n5775_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4115),
    .Q_t(n4115_t)
  );


  nnd2s3
  U2787
  (
    .DIN1(n4118),
    .DIN1_t(n4118_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4113),
    .Q_t(n4113_t)
  );


  nnd2s3
  U2788
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2166),
    .DIN2_t(n2166_t),
    .Q(n4112),
    .Q_t(n4112_t)
  );


  nnd2s3
  U2789
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2123),
    .DIN2_t(n2123_t),
    .Q(n4111),
    .Q_t(n4111_t)
  );


  nnd4s2
  U2790
  (
    .DIN1(n4119),
    .DIN1_t(n4119_t),
    .DIN2(n4120),
    .DIN2_t(n4120_t),
    .DIN3(n4121),
    .DIN3_t(n4121_t),
    .DIN4(n4122),
    .DIN4_t(n4122_t),
    .Q(WX3248),
    .Q_t(WX3248_t)
  );


  nnd2s3
  U2791
  (
    .DIN1(n3851),
    .DIN1_t(n3851_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4122),
    .Q_t(n4122_t)
  );


  xor2s3
  U2792
  (
    .DIN1(n4123),
    .DIN1_t(n4123_t),
    .DIN2(n4124),
    .DIN2_t(n4124_t),
    .Q(n3851),
    .Q_t(n3851_t)
  );


  xor2s3
  U2793
  (
    .DIN1(n5779),
    .DIN1_t(n5779_t),
    .DIN2(n4125),
    .DIN2_t(n4125_t),
    .Q(n4124),
    .Q_t(n4124_t)
  );


  xor2s3
  U2794
  (
    .DIN1(n5777),
    .DIN1_t(n5777_t),
    .DIN2(n5778),
    .DIN2_t(n5778_t),
    .Q(n4125),
    .Q_t(n4125_t)
  );


  xor2s3
  U2795
  (
    .DIN1(n5780),
    .DIN1_t(n5780_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4123),
    .Q_t(n4123_t)
  );


  nnd2s3
  U2796
  (
    .DIN1(n4126),
    .DIN1_t(n4126_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4121),
    .Q_t(n4121_t)
  );


  nnd2s3
  U2797
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2167),
    .DIN2_t(n2167_t),
    .Q(n4120),
    .Q_t(n4120_t)
  );


  nnd2s3
  U2798
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2122),
    .DIN2_t(n2122_t),
    .Q(n4119),
    .Q_t(n4119_t)
  );


  nnd4s2
  U2799
  (
    .DIN1(n4127),
    .DIN1_t(n4127_t),
    .DIN2(n4128),
    .DIN2_t(n4128_t),
    .DIN3(n4129),
    .DIN3_t(n4129_t),
    .DIN4(n4130),
    .DIN4_t(n4130_t),
    .Q(WX3246),
    .Q_t(WX3246_t)
  );


  nnd2s3
  U2800
  (
    .DIN1(n3859),
    .DIN1_t(n3859_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4130),
    .Q_t(n4130_t)
  );


  xor2s3
  U2801
  (
    .DIN1(n4131),
    .DIN1_t(n4131_t),
    .DIN2(n4132),
    .DIN2_t(n4132_t),
    .Q(n3859),
    .Q_t(n3859_t)
  );


  xor2s3
  U2802
  (
    .DIN1(n5784),
    .DIN1_t(n5784_t),
    .DIN2(n4133),
    .DIN2_t(n4133_t),
    .Q(n4132),
    .Q_t(n4132_t)
  );


  xor2s3
  U2803
  (
    .DIN1(n5782),
    .DIN1_t(n5782_t),
    .DIN2(n5783),
    .DIN2_t(n5783_t),
    .Q(n4133),
    .Q_t(n4133_t)
  );


  xor2s3
  U2804
  (
    .DIN1(n5785),
    .DIN1_t(n5785_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4131),
    .Q_t(n4131_t)
  );


  nnd2s3
  U2805
  (
    .DIN1(n4134),
    .DIN1_t(n4134_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4129),
    .Q_t(n4129_t)
  );


  nnd2s3
  U2806
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2168),
    .DIN2_t(n2168_t),
    .Q(n4128),
    .Q_t(n4128_t)
  );


  nnd2s3
  U2807
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2121),
    .DIN2_t(n2121_t),
    .Q(n4127),
    .Q_t(n4127_t)
  );


  nnd4s2
  U2808
  (
    .DIN1(n4135),
    .DIN1_t(n4135_t),
    .DIN2(n4136),
    .DIN2_t(n4136_t),
    .DIN3(n4137),
    .DIN3_t(n4137_t),
    .DIN4(n4138),
    .DIN4_t(n4138_t),
    .Q(WX3244),
    .Q_t(WX3244_t)
  );


  nnd2s3
  U2809
  (
    .DIN1(n3867),
    .DIN1_t(n3867_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4138),
    .Q_t(n4138_t)
  );


  xor2s3
  U2810
  (
    .DIN1(n4139),
    .DIN1_t(n4139_t),
    .DIN2(n4140),
    .DIN2_t(n4140_t),
    .Q(n3867),
    .Q_t(n3867_t)
  );


  xor2s3
  U2811
  (
    .DIN1(n5789),
    .DIN1_t(n5789_t),
    .DIN2(n4141),
    .DIN2_t(n4141_t),
    .Q(n4140),
    .Q_t(n4140_t)
  );


  xor2s3
  U2812
  (
    .DIN1(n5787),
    .DIN1_t(n5787_t),
    .DIN2(n5788),
    .DIN2_t(n5788_t),
    .Q(n4141),
    .Q_t(n4141_t)
  );


  xor2s3
  U2813
  (
    .DIN1(n5790),
    .DIN1_t(n5790_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4139),
    .Q_t(n4139_t)
  );


  nnd2s3
  U2814
  (
    .DIN1(n4142),
    .DIN1_t(n4142_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4137),
    .Q_t(n4137_t)
  );


  nnd2s3
  U2815
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2169),
    .DIN2_t(n2169_t),
    .Q(n4136),
    .Q_t(n4136_t)
  );


  nnd2s3
  U2816
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2120),
    .DIN2_t(n2120_t),
    .Q(n4135),
    .Q_t(n4135_t)
  );


  nnd4s2
  U2817
  (
    .DIN1(n4143),
    .DIN1_t(n4143_t),
    .DIN2(n4144),
    .DIN2_t(n4144_t),
    .DIN3(n4145),
    .DIN3_t(n4145_t),
    .DIN4(n4146),
    .DIN4_t(n4146_t),
    .Q(WX3242),
    .Q_t(WX3242_t)
  );


  nnd2s3
  U2818
  (
    .DIN1(n3875),
    .DIN1_t(n3875_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4146),
    .Q_t(n4146_t)
  );


  xor2s3
  U2819
  (
    .DIN1(n4147),
    .DIN1_t(n4147_t),
    .DIN2(n4148),
    .DIN2_t(n4148_t),
    .Q(n3875),
    .Q_t(n3875_t)
  );


  xor2s3
  U2820
  (
    .DIN1(n5794),
    .DIN1_t(n5794_t),
    .DIN2(n4149),
    .DIN2_t(n4149_t),
    .Q(n4148),
    .Q_t(n4148_t)
  );


  xor2s3
  U2821
  (
    .DIN1(n5792),
    .DIN1_t(n5792_t),
    .DIN2(n5793),
    .DIN2_t(n5793_t),
    .Q(n4149),
    .Q_t(n4149_t)
  );


  xor2s3
  U2822
  (
    .DIN1(n5795),
    .DIN1_t(n5795_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4147),
    .Q_t(n4147_t)
  );


  nnd2s3
  U2823
  (
    .DIN1(n4150),
    .DIN1_t(n4150_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4145),
    .Q_t(n4145_t)
  );


  nnd2s3
  U2824
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2170),
    .DIN2_t(n2170_t),
    .Q(n4144),
    .Q_t(n4144_t)
  );


  nnd2s3
  U2825
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2119),
    .DIN2_t(n2119_t),
    .Q(n4143),
    .Q_t(n4143_t)
  );


  nnd4s2
  U2826
  (
    .DIN1(n4151),
    .DIN1_t(n4151_t),
    .DIN2(n4152),
    .DIN2_t(n4152_t),
    .DIN3(n4153),
    .DIN3_t(n4153_t),
    .DIN4(n4154),
    .DIN4_t(n4154_t),
    .Q(WX3240),
    .Q_t(WX3240_t)
  );


  nnd2s3
  U2827
  (
    .DIN1(n3883),
    .DIN1_t(n3883_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4154),
    .Q_t(n4154_t)
  );


  xor2s3
  U2828
  (
    .DIN1(n4155),
    .DIN1_t(n4155_t),
    .DIN2(n4156),
    .DIN2_t(n4156_t),
    .Q(n3883),
    .Q_t(n3883_t)
  );


  xor2s3
  U2829
  (
    .DIN1(n5799),
    .DIN1_t(n5799_t),
    .DIN2(n4157),
    .DIN2_t(n4157_t),
    .Q(n4156),
    .Q_t(n4156_t)
  );


  xor2s3
  U2830
  (
    .DIN1(n5797),
    .DIN1_t(n5797_t),
    .DIN2(n5798),
    .DIN2_t(n5798_t),
    .Q(n4157),
    .Q_t(n4157_t)
  );


  xor2s3
  U2831
  (
    .DIN1(n5800),
    .DIN1_t(n5800_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4155),
    .Q_t(n4155_t)
  );


  nnd2s3
  U2832
  (
    .DIN1(n4158),
    .DIN1_t(n4158_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4153),
    .Q_t(n4153_t)
  );


  nnd2s3
  U2833
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2171),
    .DIN2_t(n2171_t),
    .Q(n4152),
    .Q_t(n4152_t)
  );


  nnd2s3
  U2834
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2118),
    .DIN2_t(n2118_t),
    .Q(n4151),
    .Q_t(n4151_t)
  );


  nnd4s2
  U2835
  (
    .DIN1(n4159),
    .DIN1_t(n4159_t),
    .DIN2(n4160),
    .DIN2_t(n4160_t),
    .DIN3(n4161),
    .DIN3_t(n4161_t),
    .DIN4(n4162),
    .DIN4_t(n4162_t),
    .Q(WX3238),
    .Q_t(WX3238_t)
  );


  nnd2s3
  U2836
  (
    .DIN1(n3891),
    .DIN1_t(n3891_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4162),
    .Q_t(n4162_t)
  );


  xor2s3
  U2837
  (
    .DIN1(n4163),
    .DIN1_t(n4163_t),
    .DIN2(n4164),
    .DIN2_t(n4164_t),
    .Q(n3891),
    .Q_t(n3891_t)
  );


  xor2s3
  U2838
  (
    .DIN1(n5804),
    .DIN1_t(n5804_t),
    .DIN2(n4165),
    .DIN2_t(n4165_t),
    .Q(n4164),
    .Q_t(n4164_t)
  );


  xor2s3
  U2839
  (
    .DIN1(n5802),
    .DIN1_t(n5802_t),
    .DIN2(n5803),
    .DIN2_t(n5803_t),
    .Q(n4165),
    .Q_t(n4165_t)
  );


  xor2s3
  U2840
  (
    .DIN1(n5805),
    .DIN1_t(n5805_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4163),
    .Q_t(n4163_t)
  );


  nnd2s3
  U2841
  (
    .DIN1(n4166),
    .DIN1_t(n4166_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4161),
    .Q_t(n4161_t)
  );


  nnd2s3
  U2842
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2172),
    .DIN2_t(n2172_t),
    .Q(n4160),
    .Q_t(n4160_t)
  );


  nnd2s3
  U2843
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2117),
    .DIN2_t(n2117_t),
    .Q(n4159),
    .Q_t(n4159_t)
  );


  nnd4s2
  U2844
  (
    .DIN1(n4167),
    .DIN1_t(n4167_t),
    .DIN2(n4168),
    .DIN2_t(n4168_t),
    .DIN3(n4169),
    .DIN3_t(n4169_t),
    .DIN4(n4170),
    .DIN4_t(n4170_t),
    .Q(WX3236),
    .Q_t(WX3236_t)
  );


  nnd2s3
  U2845
  (
    .DIN1(n3899),
    .DIN1_t(n3899_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4170),
    .Q_t(n4170_t)
  );


  xor2s3
  U2846
  (
    .DIN1(n4171),
    .DIN1_t(n4171_t),
    .DIN2(n4172),
    .DIN2_t(n4172_t),
    .Q(n3899),
    .Q_t(n3899_t)
  );


  xor2s3
  U2847
  (
    .DIN1(n5809),
    .DIN1_t(n5809_t),
    .DIN2(n4173),
    .DIN2_t(n4173_t),
    .Q(n4172),
    .Q_t(n4172_t)
  );


  xor2s3
  U2848
  (
    .DIN1(n5807),
    .DIN1_t(n5807_t),
    .DIN2(n5808),
    .DIN2_t(n5808_t),
    .Q(n4173),
    .Q_t(n4173_t)
  );


  xor2s3
  U2849
  (
    .DIN1(n5810),
    .DIN1_t(n5810_t),
    .DIN2(n6692),
    .DIN2_t(n6692_t),
    .Q(n4171),
    .Q_t(n4171_t)
  );


  nnd2s3
  U2850
  (
    .DIN1(n4174),
    .DIN1_t(n4174_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4169),
    .Q_t(n4169_t)
  );


  nnd2s3
  U2851
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2173),
    .DIN2_t(n2173_t),
    .Q(n4168),
    .Q_t(n4168_t)
  );


  nnd2s3
  U2852
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2116),
    .DIN2_t(n2116_t),
    .Q(n4167),
    .Q_t(n4167_t)
  );


  nnd4s2
  U2853
  (
    .DIN1(n4175),
    .DIN1_t(n4175_t),
    .DIN2(n4176),
    .DIN2_t(n4176_t),
    .DIN3(n4177),
    .DIN3_t(n4177_t),
    .DIN4(n4178),
    .DIN4_t(n4178_t),
    .Q(WX3234),
    .Q_t(WX3234_t)
  );


  nnd2s3
  U2854
  (
    .DIN1(n3907),
    .DIN1_t(n3907_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4178),
    .Q_t(n4178_t)
  );


  xor2s3
  U2855
  (
    .DIN1(n4179),
    .DIN1_t(n4179_t),
    .DIN2(n4180),
    .DIN2_t(n4180_t),
    .Q(n3907),
    .Q_t(n3907_t)
  );


  xor2s3
  U2856
  (
    .DIN1(n5814),
    .DIN1_t(n5814_t),
    .DIN2(n4181),
    .DIN2_t(n4181_t),
    .Q(n4180),
    .Q_t(n4180_t)
  );


  xor2s3
  U2857
  (
    .DIN1(n5812),
    .DIN1_t(n5812_t),
    .DIN2(n5813),
    .DIN2_t(n5813_t),
    .Q(n4181),
    .Q_t(n4181_t)
  );


  xor2s3
  U2858
  (
    .DIN1(n5815),
    .DIN1_t(n5815_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4179),
    .Q_t(n4179_t)
  );


  nnd2s3
  U2859
  (
    .DIN1(n4182),
    .DIN1_t(n4182_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4177),
    .Q_t(n4177_t)
  );


  nnd2s3
  U2860
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2174),
    .DIN2_t(n2174_t),
    .Q(n4176),
    .Q_t(n4176_t)
  );


  nnd2s3
  U2861
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2115),
    .DIN2_t(n2115_t),
    .Q(n4175),
    .Q_t(n4175_t)
  );


  nnd4s2
  U2862
  (
    .DIN1(n4183),
    .DIN1_t(n4183_t),
    .DIN2(n4184),
    .DIN2_t(n4184_t),
    .DIN3(n4185),
    .DIN3_t(n4185_t),
    .DIN4(n4186),
    .DIN4_t(n4186_t),
    .Q(WX3232),
    .Q_t(WX3232_t)
  );


  nnd2s3
  U2863
  (
    .DIN1(n3915),
    .DIN1_t(n3915_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4186),
    .Q_t(n4186_t)
  );


  xor2s3
  U2864
  (
    .DIN1(n4187),
    .DIN1_t(n4187_t),
    .DIN2(n4188),
    .DIN2_t(n4188_t),
    .Q(n3915),
    .Q_t(n3915_t)
  );


  xor2s3
  U2865
  (
    .DIN1(n5819),
    .DIN1_t(n5819_t),
    .DIN2(n4189),
    .DIN2_t(n4189_t),
    .Q(n4188),
    .Q_t(n4188_t)
  );


  xor2s3
  U2866
  (
    .DIN1(n5817),
    .DIN1_t(n5817_t),
    .DIN2(n5818),
    .DIN2_t(n5818_t),
    .Q(n4189),
    .Q_t(n4189_t)
  );


  xor2s3
  U2867
  (
    .DIN1(n5820),
    .DIN1_t(n5820_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4187),
    .Q_t(n4187_t)
  );


  nnd2s3
  U2868
  (
    .DIN1(n4190),
    .DIN1_t(n4190_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4185),
    .Q_t(n4185_t)
  );


  nnd2s3
  U2869
  (
    .DIN1(n6599),
    .DIN1_t(n6599_t),
    .DIN2(n2175),
    .DIN2_t(n2175_t),
    .Q(n4184),
    .Q_t(n4184_t)
  );


  nnd2s3
  U2870
  (
    .DIN1(n6568),
    .DIN1_t(n6568_t),
    .DIN2(n2114),
    .DIN2_t(n2114_t),
    .Q(n4183),
    .Q_t(n4183_t)
  );


  nnd4s2
  U2871
  (
    .DIN1(n4191),
    .DIN1_t(n4191_t),
    .DIN2(n4192),
    .DIN2_t(n4192_t),
    .DIN3(n4193),
    .DIN3_t(n4193_t),
    .DIN4(n4194),
    .DIN4_t(n4194_t),
    .Q(WX3230),
    .Q_t(WX3230_t)
  );


  nnd2s3
  U2872
  (
    .DIN1(n3923),
    .DIN1_t(n3923_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4194),
    .Q_t(n4194_t)
  );


  xor2s3
  U2873
  (
    .DIN1(n4195),
    .DIN1_t(n4195_t),
    .DIN2(n4196),
    .DIN2_t(n4196_t),
    .Q(n3923),
    .Q_t(n3923_t)
  );


  xor2s3
  U2874
  (
    .DIN1(n5824),
    .DIN1_t(n5824_t),
    .DIN2(n4197),
    .DIN2_t(n4197_t),
    .Q(n4196),
    .Q_t(n4196_t)
  );


  xor2s3
  U2875
  (
    .DIN1(n5822),
    .DIN1_t(n5822_t),
    .DIN2(n5823),
    .DIN2_t(n5823_t),
    .Q(n4197),
    .Q_t(n4197_t)
  );


  xor2s3
  U2876
  (
    .DIN1(n5825),
    .DIN1_t(n5825_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4195),
    .Q_t(n4195_t)
  );


  nnd2s3
  U2877
  (
    .DIN1(n4198),
    .DIN1_t(n4198_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4193),
    .Q_t(n4193_t)
  );


  nnd2s3
  U2878
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2176),
    .DIN2_t(n2176_t),
    .Q(n4192),
    .Q_t(n4192_t)
  );


  nnd2s3
  U2879
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2113),
    .DIN2_t(n2113_t),
    .Q(n4191),
    .Q_t(n4191_t)
  );


  nor2s3
  U2880
  (
    .DIN1(n6802),
    .DIN1_t(n6802_t),
    .DIN2(n2176),
    .DIN2_t(n2176_t),
    .Q(WX3132),
    .Q_t(WX3132_t)
  );


  nor2s3
  U2881
  (
    .DIN1(n5828),
    .DIN1_t(n5828_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3130),
    .Q_t(WX3130_t)
  );


  nor2s3
  U2882
  (
    .DIN1(n5829),
    .DIN1_t(n5829_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3128),
    .Q_t(WX3128_t)
  );


  nor2s3
  U2883
  (
    .DIN1(n5830),
    .DIN1_t(n5830_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3126),
    .Q_t(WX3126_t)
  );


  nor2s3
  U2884
  (
    .DIN1(n5831),
    .DIN1_t(n5831_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3124),
    .Q_t(WX3124_t)
  );


  nor2s3
  U2885
  (
    .DIN1(n5832),
    .DIN1_t(n5832_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3122),
    .Q_t(WX3122_t)
  );


  nor2s3
  U2886
  (
    .DIN1(n5833),
    .DIN1_t(n5833_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3120),
    .Q_t(WX3120_t)
  );


  nor2s3
  U2887
  (
    .DIN1(n5834),
    .DIN1_t(n5834_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3118),
    .Q_t(WX3118_t)
  );


  nor2s3
  U2888
  (
    .DIN1(n5835),
    .DIN1_t(n5835_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3116),
    .Q_t(WX3116_t)
  );


  nor2s3
  U2889
  (
    .DIN1(n5836),
    .DIN1_t(n5836_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3114),
    .Q_t(WX3114_t)
  );


  nor2s3
  U2890
  (
    .DIN1(n5837),
    .DIN1_t(n5837_t),
    .DIN2(n6765),
    .DIN2_t(n6765_t),
    .Q(WX3112),
    .Q_t(WX3112_t)
  );


  nor2s3
  U2891
  (
    .DIN1(n5838),
    .DIN1_t(n5838_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3110),
    .Q_t(WX3110_t)
  );


  nor2s3
  U2892
  (
    .DIN1(n5839),
    .DIN1_t(n5839_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3108),
    .Q_t(WX3108_t)
  );


  nor2s3
  U2893
  (
    .DIN1(n5840),
    .DIN1_t(n5840_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3106),
    .Q_t(WX3106_t)
  );


  nor2s3
  U2894
  (
    .DIN1(n5841),
    .DIN1_t(n5841_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3104),
    .Q_t(WX3104_t)
  );


  nor2s3
  U2895
  (
    .DIN1(n5842),
    .DIN1_t(n5842_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3102),
    .Q_t(WX3102_t)
  );


  nor2s3
  U2896
  (
    .DIN1(n5843),
    .DIN1_t(n5843_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3100),
    .Q_t(WX3100_t)
  );


  nor2s3
  U2897
  (
    .DIN1(n5844),
    .DIN1_t(n5844_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3098),
    .Q_t(WX3098_t)
  );


  nor2s3
  U2898
  (
    .DIN1(n5845),
    .DIN1_t(n5845_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3096),
    .Q_t(WX3096_t)
  );


  nor2s3
  U2899
  (
    .DIN1(n5846),
    .DIN1_t(n5846_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3094),
    .Q_t(WX3094_t)
  );


  nor2s3
  U2900
  (
    .DIN1(n5847),
    .DIN1_t(n5847_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3092),
    .Q_t(WX3092_t)
  );


  nor2s3
  U2901
  (
    .DIN1(n5848),
    .DIN1_t(n5848_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3090),
    .Q_t(WX3090_t)
  );


  nor2s3
  U2902
  (
    .DIN1(n5849),
    .DIN1_t(n5849_t),
    .DIN2(n6764),
    .DIN2_t(n6764_t),
    .Q(WX3088),
    .Q_t(WX3088_t)
  );


  nor2s3
  U2903
  (
    .DIN1(n5850),
    .DIN1_t(n5850_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX3086),
    .Q_t(WX3086_t)
  );


  nor2s3
  U2904
  (
    .DIN1(n5851),
    .DIN1_t(n5851_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX3084),
    .Q_t(WX3084_t)
  );


  nor2s3
  U2905
  (
    .DIN1(n5852),
    .DIN1_t(n5852_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX3082),
    .Q_t(WX3082_t)
  );


  nor2s3
  U2906
  (
    .DIN1(n5853),
    .DIN1_t(n5853_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX3080),
    .Q_t(WX3080_t)
  );


  nor2s3
  U2907
  (
    .DIN1(n5854),
    .DIN1_t(n5854_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX3078),
    .Q_t(WX3078_t)
  );


  nor2s3
  U2908
  (
    .DIN1(n5855),
    .DIN1_t(n5855_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX3076),
    .Q_t(WX3076_t)
  );


  nor2s3
  U2909
  (
    .DIN1(n5856),
    .DIN1_t(n5856_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX3074),
    .Q_t(WX3074_t)
  );


  nor2s3
  U2910
  (
    .DIN1(n5857),
    .DIN1_t(n5857_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX3072),
    .Q_t(WX3072_t)
  );


  nor2s3
  U2911
  (
    .DIN1(n5858),
    .DIN1_t(n5858_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX3070),
    .Q_t(WX3070_t)
  );


  nor2s3
  U2912
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n4199),
    .DIN2_t(n4199_t),
    .Q(WX2619),
    .Q_t(WX2619_t)
  );


  xor2s3
  U2913
  (
    .DIN1(n6105),
    .DIN1_t(n6105_t),
    .DIN2(n6113),
    .DIN2_t(n6113_t),
    .Q(n4199),
    .Q_t(n4199_t)
  );


  nor2s3
  U2914
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n4200),
    .DIN2_t(n4200_t),
    .Q(WX2617),
    .Q_t(WX2617_t)
  );


  xor2s3
  U2915
  (
    .DIN1(n6096),
    .DIN1_t(n6096_t),
    .DIN2(n6104),
    .DIN2_t(n6104_t),
    .Q(n4200),
    .Q_t(n4200_t)
  );


  nor2s3
  U2916
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n4201),
    .DIN2_t(n4201_t),
    .Q(WX2615),
    .Q_t(WX2615_t)
  );


  xor2s3
  U2917
  (
    .DIN1(n6087),
    .DIN1_t(n6087_t),
    .DIN2(n6095),
    .DIN2_t(n6095_t),
    .Q(n4201),
    .Q_t(n4201_t)
  );


  nor2s3
  U2918
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n4202),
    .DIN2_t(n4202_t),
    .Q(WX2613),
    .Q_t(WX2613_t)
  );


  xor2s3
  U2919
  (
    .DIN1(n6078),
    .DIN1_t(n6078_t),
    .DIN2(n6086),
    .DIN2_t(n6086_t),
    .Q(n4202),
    .Q_t(n4202_t)
  );


  nor2s3
  U2920
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n4203),
    .DIN2_t(n4203_t),
    .Q(WX2611),
    .Q_t(WX2611_t)
  );


  xor2s3
  U2921
  (
    .DIN1(n6069),
    .DIN1_t(n6069_t),
    .DIN2(n6077),
    .DIN2_t(n6077_t),
    .Q(n4203),
    .Q_t(n4203_t)
  );


  nor2s3
  U2922
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n4204),
    .DIN2_t(n4204_t),
    .Q(WX2609),
    .Q_t(WX2609_t)
  );


  xor2s3
  U2923
  (
    .DIN1(n6060),
    .DIN1_t(n6060_t),
    .DIN2(n6068),
    .DIN2_t(n6068_t),
    .Q(n4204),
    .Q_t(n4204_t)
  );


  nor2s3
  U2924
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n4205),
    .DIN2_t(n4205_t),
    .Q(WX2607),
    .Q_t(WX2607_t)
  );


  xor2s3
  U2925
  (
    .DIN1(n6051),
    .DIN1_t(n6051_t),
    .DIN2(n6059),
    .DIN2_t(n6059_t),
    .Q(n4205),
    .Q_t(n4205_t)
  );


  nor2s3
  U2926
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n4206),
    .DIN2_t(n4206_t),
    .Q(WX2605),
    .Q_t(WX2605_t)
  );


  xor2s3
  U2927
  (
    .DIN1(n6042),
    .DIN1_t(n6042_t),
    .DIN2(n6050),
    .DIN2_t(n6050_t),
    .Q(n4206),
    .Q_t(n4206_t)
  );


  nor2s3
  U2928
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n4207),
    .DIN2_t(n4207_t),
    .Q(WX2603),
    .Q_t(WX2603_t)
  );


  xor2s3
  U2929
  (
    .DIN1(n6033),
    .DIN1_t(n6033_t),
    .DIN2(n6041),
    .DIN2_t(n6041_t),
    .Q(n4207),
    .Q_t(n4207_t)
  );


  nor2s3
  U2930
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n4208),
    .DIN2_t(n4208_t),
    .Q(WX2601),
    .Q_t(WX2601_t)
  );


  xor2s3
  U2931
  (
    .DIN1(n6024),
    .DIN1_t(n6024_t),
    .DIN2(n6032),
    .DIN2_t(n6032_t),
    .Q(n4208),
    .Q_t(n4208_t)
  );


  nor2s3
  U2932
  (
    .DIN1(n6796),
    .DIN1_t(n6796_t),
    .DIN2(n4209),
    .DIN2_t(n4209_t),
    .Q(WX2599),
    .Q_t(WX2599_t)
  );


  xor2s3
  U2933
  (
    .DIN1(n6015),
    .DIN1_t(n6015_t),
    .DIN2(n6023),
    .DIN2_t(n6023_t),
    .Q(n4209),
    .Q_t(n4209_t)
  );


  nor2s3
  U2934
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n4210),
    .DIN2_t(n4210_t),
    .Q(WX2597),
    .Q_t(WX2597_t)
  );


  xor2s3
  U2935
  (
    .DIN1(n6006),
    .DIN1_t(n6006_t),
    .DIN2(n6014),
    .DIN2_t(n6014_t),
    .Q(n4210),
    .Q_t(n4210_t)
  );


  nor2s3
  U2936
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n4211),
    .DIN2_t(n4211_t),
    .Q(WX2595),
    .Q_t(WX2595_t)
  );


  xor2s3
  U2937
  (
    .DIN1(n5997),
    .DIN1_t(n5997_t),
    .DIN2(n6005),
    .DIN2_t(n6005_t),
    .Q(n4211),
    .Q_t(n4211_t)
  );


  nor2s3
  U2938
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n4212),
    .DIN2_t(n4212_t),
    .Q(WX2593),
    .Q_t(WX2593_t)
  );


  xor2s3
  U2939
  (
    .DIN1(n5988),
    .DIN1_t(n5988_t),
    .DIN2(n5996),
    .DIN2_t(n5996_t),
    .Q(n4212),
    .Q_t(n4212_t)
  );


  nor2s3
  U2940
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n4213),
    .DIN2_t(n4213_t),
    .Q(WX2591),
    .Q_t(WX2591_t)
  );


  xor2s3
  U2941
  (
    .DIN1(n5979),
    .DIN1_t(n5979_t),
    .DIN2(n5987),
    .DIN2_t(n5987_t),
    .Q(n4213),
    .Q_t(n4213_t)
  );


  nor2s3
  U2942
  (
    .DIN1(n4214),
    .DIN1_t(n4214_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX2589),
    .Q_t(WX2589_t)
  );


  xor2s3
  U2943
  (
    .DIN1(n2177),
    .DIN1_t(n2177_t),
    .DIN2(n4215),
    .DIN2_t(n4215_t),
    .Q(n4214),
    .Q_t(n4214_t)
  );


  xor2s3
  U2944
  (
    .DIN1(n5970),
    .DIN1_t(n5970_t),
    .DIN2(n5978),
    .DIN2_t(n5978_t),
    .Q(n4215),
    .Q_t(n4215_t)
  );


  nor2s3
  U2945
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n4216),
    .DIN2_t(n4216_t),
    .Q(WX2587),
    .Q_t(WX2587_t)
  );


  xor2s3
  U2946
  (
    .DIN1(n5963),
    .DIN1_t(n5963_t),
    .DIN2(n3316),
    .DIN2_t(n3316_t),
    .Q(n4216),
    .Q_t(n4216_t)
  );


  nor2s3
  U2947
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n4217),
    .DIN2_t(n4217_t),
    .Q(WX2585),
    .Q_t(WX2585_t)
  );


  xor2s3
  U2948
  (
    .DIN1(n5956),
    .DIN1_t(n5956_t),
    .DIN2(n3314),
    .DIN2_t(n3314_t),
    .Q(n4217),
    .Q_t(n4217_t)
  );


  nor2s3
  U2949
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n4218),
    .DIN2_t(n4218_t),
    .Q(WX2583),
    .Q_t(WX2583_t)
  );


  xor2s3
  U2950
  (
    .DIN1(n5949),
    .DIN1_t(n5949_t),
    .DIN2(n3312),
    .DIN2_t(n3312_t),
    .Q(n4218),
    .Q_t(n4218_t)
  );


  nor2s3
  U2951
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n4219),
    .DIN2_t(n4219_t),
    .Q(WX2581),
    .Q_t(WX2581_t)
  );


  xor2s3
  U2952
  (
    .DIN1(n5942),
    .DIN1_t(n5942_t),
    .DIN2(n3310),
    .DIN2_t(n3310_t),
    .Q(n4219),
    .Q_t(n4219_t)
  );


  nor2s3
  U2953
  (
    .DIN1(n4220),
    .DIN1_t(n4220_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX2579),
    .Q_t(WX2579_t)
  );


  xnr2s3
  U2954
  (
    .DIN1(n3308),
    .DIN1_t(n3308_t),
    .DIN2(n4221),
    .DIN2_t(n4221_t),
    .Q(n4220),
    .Q_t(n4220_t)
  );


  xor2s3
  U2955
  (
    .DIN1(n5935),
    .DIN1_t(n5935_t),
    .DIN2(n6114),
    .DIN2_t(n6114_t),
    .Q(n4221),
    .Q_t(n4221_t)
  );


  nor2s3
  U2956
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n4222),
    .DIN2_t(n4222_t),
    .Q(WX2577),
    .Q_t(WX2577_t)
  );


  xor2s3
  U2957
  (
    .DIN1(n5928),
    .DIN1_t(n5928_t),
    .DIN2(n3306),
    .DIN2_t(n3306_t),
    .Q(n4222),
    .Q_t(n4222_t)
  );


  nor2s3
  U2958
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n4223),
    .DIN2_t(n4223_t),
    .Q(WX2575),
    .Q_t(WX2575_t)
  );


  xor2s3
  U2959
  (
    .DIN1(n5921),
    .DIN1_t(n5921_t),
    .DIN2(n3304),
    .DIN2_t(n3304_t),
    .Q(n4223),
    .Q_t(n4223_t)
  );


  nor2s3
  U2960
  (
    .DIN1(n6797),
    .DIN1_t(n6797_t),
    .DIN2(n4224),
    .DIN2_t(n4224_t),
    .Q(WX2573),
    .Q_t(WX2573_t)
  );


  xor2s3
  U2961
  (
    .DIN1(n5914),
    .DIN1_t(n5914_t),
    .DIN2(n3302),
    .DIN2_t(n3302_t),
    .Q(n4224),
    .Q_t(n4224_t)
  );


  nor2s3
  U2962
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n4225),
    .DIN2_t(n4225_t),
    .Q(WX2571),
    .Q_t(WX2571_t)
  );


  xor2s3
  U2963
  (
    .DIN1(n5907),
    .DIN1_t(n5907_t),
    .DIN2(n3300),
    .DIN2_t(n3300_t),
    .Q(n4225),
    .Q_t(n4225_t)
  );


  nor2s3
  U2964
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n4226),
    .DIN2_t(n4226_t),
    .Q(WX2569),
    .Q_t(WX2569_t)
  );


  xor2s3
  U2965
  (
    .DIN1(n5900),
    .DIN1_t(n5900_t),
    .DIN2(n3298),
    .DIN2_t(n3298_t),
    .Q(n4226),
    .Q_t(n4226_t)
  );


  nor2s3
  U2966
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n4227),
    .DIN2_t(n4227_t),
    .Q(WX2567),
    .Q_t(WX2567_t)
  );


  xor2s3
  U2967
  (
    .DIN1(n5893),
    .DIN1_t(n5893_t),
    .DIN2(n3296),
    .DIN2_t(n3296_t),
    .Q(n4227),
    .Q_t(n4227_t)
  );


  nor2s3
  U2968
  (
    .DIN1(n4228),
    .DIN1_t(n4228_t),
    .DIN2(n6763),
    .DIN2_t(n6763_t),
    .Q(WX2565),
    .Q_t(WX2565_t)
  );


  xnr2s3
  U2969
  (
    .DIN1(n3294),
    .DIN1_t(n3294_t),
    .DIN2(n4229),
    .DIN2_t(n4229_t),
    .Q(n4228),
    .Q_t(n4228_t)
  );


  xor2s3
  U2970
  (
    .DIN1(n5886),
    .DIN1_t(n5886_t),
    .DIN2(n6114),
    .DIN2_t(n6114_t),
    .Q(n4229),
    .Q_t(n4229_t)
  );


  nor2s3
  U2971
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n4230),
    .DIN2_t(n4230_t),
    .Q(WX2563),
    .Q_t(WX2563_t)
  );


  xor2s3
  U2972
  (
    .DIN1(n5879),
    .DIN1_t(n5879_t),
    .DIN2(n3292),
    .DIN2_t(n3292_t),
    .Q(n4230),
    .Q_t(n4230_t)
  );


  nor2s3
  U2973
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n4231),
    .DIN2_t(n4231_t),
    .Q(WX2561),
    .Q_t(WX2561_t)
  );


  xor2s3
  U2974
  (
    .DIN1(n5872),
    .DIN1_t(n5872_t),
    .DIN2(n3290),
    .DIN2_t(n3290_t),
    .Q(n4231),
    .Q_t(n4231_t)
  );


  nor2s3
  U2975
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n4232),
    .DIN2_t(n4232_t),
    .Q(WX2559),
    .Q_t(WX2559_t)
  );


  xor2s3
  U2976
  (
    .DIN1(n5865),
    .DIN1_t(n5865_t),
    .DIN2(n3288),
    .DIN2_t(n3288_t),
    .Q(n4232),
    .Q_t(n4232_t)
  );


  nor2s3
  U2977
  (
    .DIN1(n6798),
    .DIN1_t(n6798_t),
    .DIN2(n4233),
    .DIN2_t(n4233_t),
    .Q(WX2557),
    .Q_t(WX2557_t)
  );


  xor2s3
  U2978
  (
    .DIN1(n6114),
    .DIN1_t(n6114_t),
    .DIN2(n3286),
    .DIN2_t(n3286_t),
    .Q(n4233),
    .Q_t(n4233_t)
  );


  nor2s3
  U2979
  (
    .DIN1(n5864),
    .DIN1_t(n5864_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2191),
    .Q_t(WX2191_t)
  );


  nor2s3
  U2980
  (
    .DIN1(n5871),
    .DIN1_t(n5871_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2189),
    .Q_t(WX2189_t)
  );


  nor2s3
  U2981
  (
    .DIN1(n5878),
    .DIN1_t(n5878_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2187),
    .Q_t(WX2187_t)
  );


  nor2s3
  U2982
  (
    .DIN1(n5885),
    .DIN1_t(n5885_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2185),
    .Q_t(WX2185_t)
  );


  nor2s3
  U2983
  (
    .DIN1(n5892),
    .DIN1_t(n5892_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2183),
    .Q_t(WX2183_t)
  );


  nor2s3
  U2984
  (
    .DIN1(n5899),
    .DIN1_t(n5899_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2181),
    .Q_t(WX2181_t)
  );


  nor2s3
  U2985
  (
    .DIN1(n5906),
    .DIN1_t(n5906_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2179),
    .Q_t(WX2179_t)
  );


  nor2s3
  U2986
  (
    .DIN1(n5913),
    .DIN1_t(n5913_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2177),
    .Q_t(WX2177_t)
  );


  nor2s3
  U2987
  (
    .DIN1(n5920),
    .DIN1_t(n5920_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2175),
    .Q_t(WX2175_t)
  );


  nor2s3
  U2988
  (
    .DIN1(n5927),
    .DIN1_t(n5927_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2173),
    .Q_t(WX2173_t)
  );


  nor2s3
  U2989
  (
    .DIN1(n5934),
    .DIN1_t(n5934_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2171),
    .Q_t(WX2171_t)
  );


  nor2s3
  U2990
  (
    .DIN1(n5941),
    .DIN1_t(n5941_t),
    .DIN2(n6762),
    .DIN2_t(n6762_t),
    .Q(WX2169),
    .Q_t(WX2169_t)
  );


  nor2s3
  U2991
  (
    .DIN1(n5948),
    .DIN1_t(n5948_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX2167),
    .Q_t(WX2167_t)
  );


  nor2s3
  U2992
  (
    .DIN1(n5955),
    .DIN1_t(n5955_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX2165),
    .Q_t(WX2165_t)
  );


  nor2s3
  U2993
  (
    .DIN1(n5962),
    .DIN1_t(n5962_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX2163),
    .Q_t(WX2163_t)
  );


  nor2s3
  U2994
  (
    .DIN1(n5969),
    .DIN1_t(n5969_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX2161),
    .Q_t(WX2161_t)
  );


  nor2s3
  U2995
  (
    .DIN1(n5977),
    .DIN1_t(n5977_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX2159),
    .Q_t(WX2159_t)
  );


  nor2s3
  U2996
  (
    .DIN1(n5986),
    .DIN1_t(n5986_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX2157),
    .Q_t(WX2157_t)
  );


  nor2s3
  U2997
  (
    .DIN1(n5995),
    .DIN1_t(n5995_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX2155),
    .Q_t(WX2155_t)
  );


  nor2s3
  U2998
  (
    .DIN1(n6004),
    .DIN1_t(n6004_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX2153),
    .Q_t(WX2153_t)
  );


  nor2s3
  U2999
  (
    .DIN1(n6013),
    .DIN1_t(n6013_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX2151),
    .Q_t(WX2151_t)
  );


  nor2s3
  U3000
  (
    .DIN1(n6022),
    .DIN1_t(n6022_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX2149),
    .Q_t(WX2149_t)
  );


  nor2s3
  U3001
  (
    .DIN1(n6031),
    .DIN1_t(n6031_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX2147),
    .Q_t(WX2147_t)
  );


  nor2s3
  U3002
  (
    .DIN1(n6040),
    .DIN1_t(n6040_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2145),
    .Q_t(WX2145_t)
  );


  nor2s3
  U3003
  (
    .DIN1(n6049),
    .DIN1_t(n6049_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2143),
    .Q_t(WX2143_t)
  );


  nor2s3
  U3004
  (
    .DIN1(n6058),
    .DIN1_t(n6058_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2141),
    .Q_t(WX2141_t)
  );


  nor2s3
  U3005
  (
    .DIN1(n6067),
    .DIN1_t(n6067_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2139),
    .Q_t(WX2139_t)
  );


  nor2s3
  U3006
  (
    .DIN1(n6076),
    .DIN1_t(n6076_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2137),
    .Q_t(WX2137_t)
  );


  nor2s3
  U3007
  (
    .DIN1(n6085),
    .DIN1_t(n6085_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2135),
    .Q_t(WX2135_t)
  );


  nor2s3
  U3008
  (
    .DIN1(n6094),
    .DIN1_t(n6094_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2133),
    .Q_t(WX2133_t)
  );


  nor2s3
  U3009
  (
    .DIN1(n6103),
    .DIN1_t(n6103_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2131),
    .Q_t(WX2131_t)
  );


  nor2s3
  U3010
  (
    .DIN1(n6112),
    .DIN1_t(n6112_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2129),
    .Q_t(WX2129_t)
  );


  and2s3
  U3011
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5863),
    .DIN2_t(n5863_t),
    .Q(WX2127),
    .Q_t(WX2127_t)
  );


  and2s3
  U3012
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5870),
    .DIN2_t(n5870_t),
    .Q(WX2125),
    .Q_t(WX2125_t)
  );


  and2s3
  U3013
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5877),
    .DIN2_t(n5877_t),
    .Q(WX2123),
    .Q_t(WX2123_t)
  );


  and2s3
  U3014
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5884),
    .DIN2_t(n5884_t),
    .Q(WX2121),
    .Q_t(WX2121_t)
  );


  and2s3
  U3015
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5891),
    .DIN2_t(n5891_t),
    .Q(WX2119),
    .Q_t(WX2119_t)
  );


  and2s3
  U3016
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5898),
    .DIN2_t(n5898_t),
    .Q(WX2117),
    .Q_t(WX2117_t)
  );


  and2s3
  U3017
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5905),
    .DIN2_t(n5905_t),
    .Q(WX2115),
    .Q_t(WX2115_t)
  );


  and2s3
  U3018
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5912),
    .DIN2_t(n5912_t),
    .Q(WX2113),
    .Q_t(WX2113_t)
  );


  and2s3
  U3019
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5919),
    .DIN2_t(n5919_t),
    .Q(WX2111),
    .Q_t(WX2111_t)
  );


  and2s3
  U3020
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5926),
    .DIN2_t(n5926_t),
    .Q(WX2109),
    .Q_t(WX2109_t)
  );


  and2s3
  U3021
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5933),
    .DIN2_t(n5933_t),
    .Q(WX2107),
    .Q_t(WX2107_t)
  );


  and2s3
  U3022
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5940),
    .DIN2_t(n5940_t),
    .Q(WX2105),
    .Q_t(WX2105_t)
  );


  and2s3
  U3023
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5947),
    .DIN2_t(n5947_t),
    .Q(WX2103),
    .Q_t(WX2103_t)
  );


  and2s3
  U3024
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5954),
    .DIN2_t(n5954_t),
    .Q(WX2101),
    .Q_t(WX2101_t)
  );


  and2s3
  U3025
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5961),
    .DIN2_t(n5961_t),
    .Q(WX2099),
    .Q_t(WX2099_t)
  );


  and2s3
  U3026
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5968),
    .DIN2_t(n5968_t),
    .Q(WX2097),
    .Q_t(WX2097_t)
  );


  and2s3
  U3027
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5976),
    .DIN2_t(n5976_t),
    .Q(WX2095),
    .Q_t(WX2095_t)
  );


  and2s3
  U3028
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5985),
    .DIN2_t(n5985_t),
    .Q(WX2093),
    .Q_t(WX2093_t)
  );


  and2s3
  U3029
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n5994),
    .DIN2_t(n5994_t),
    .Q(WX2091),
    .Q_t(WX2091_t)
  );


  and2s3
  U3030
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6003),
    .DIN2_t(n6003_t),
    .Q(WX2089),
    .Q_t(WX2089_t)
  );


  and2s3
  U3031
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6012),
    .DIN2_t(n6012_t),
    .Q(WX2087),
    .Q_t(WX2087_t)
  );


  and2s3
  U3032
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6021),
    .DIN2_t(n6021_t),
    .Q(WX2085),
    .Q_t(WX2085_t)
  );


  and2s3
  U3033
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6030),
    .DIN2_t(n6030_t),
    .Q(WX2083),
    .Q_t(WX2083_t)
  );


  and2s3
  U3034
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6039),
    .DIN2_t(n6039_t),
    .Q(WX2081),
    .Q_t(WX2081_t)
  );


  and2s3
  U3035
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6048),
    .DIN2_t(n6048_t),
    .Q(WX2079),
    .Q_t(WX2079_t)
  );


  and2s3
  U3036
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6057),
    .DIN2_t(n6057_t),
    .Q(WX2077),
    .Q_t(WX2077_t)
  );


  and2s3
  U3037
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6066),
    .DIN2_t(n6066_t),
    .Q(WX2075),
    .Q_t(WX2075_t)
  );


  and2s3
  U3038
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6075),
    .DIN2_t(n6075_t),
    .Q(WX2073),
    .Q_t(WX2073_t)
  );


  and2s3
  U3039
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6084),
    .DIN2_t(n6084_t),
    .Q(WX2071),
    .Q_t(WX2071_t)
  );


  and2s3
  U3040
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6093),
    .DIN2_t(n6093_t),
    .Q(WX2069),
    .Q_t(WX2069_t)
  );


  and2s3
  U3041
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6102),
    .DIN2_t(n6102_t),
    .Q(WX2067),
    .Q_t(WX2067_t)
  );


  and2s3
  U3042
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6111),
    .DIN2_t(n6111_t),
    .Q(WX2065),
    .Q_t(WX2065_t)
  );


  nor2s3
  U3043
  (
    .DIN1(n5862),
    .DIN1_t(n5862_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2063),
    .Q_t(WX2063_t)
  );


  nor2s3
  U3044
  (
    .DIN1(n5869),
    .DIN1_t(n5869_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2061),
    .Q_t(WX2061_t)
  );


  nor2s3
  U3045
  (
    .DIN1(n5876),
    .DIN1_t(n5876_t),
    .DIN2(n6760),
    .DIN2_t(n6760_t),
    .Q(WX2059),
    .Q_t(WX2059_t)
  );


  nor2s3
  U3046
  (
    .DIN1(n5883),
    .DIN1_t(n5883_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2057),
    .Q_t(WX2057_t)
  );


  nor2s3
  U3047
  (
    .DIN1(n5890),
    .DIN1_t(n5890_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2055),
    .Q_t(WX2055_t)
  );


  nor2s3
  U3048
  (
    .DIN1(n5897),
    .DIN1_t(n5897_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2053),
    .Q_t(WX2053_t)
  );


  nor2s3
  U3049
  (
    .DIN1(n5904),
    .DIN1_t(n5904_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2051),
    .Q_t(WX2051_t)
  );


  nor2s3
  U3050
  (
    .DIN1(n5911),
    .DIN1_t(n5911_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2049),
    .Q_t(WX2049_t)
  );


  nor2s3
  U3051
  (
    .DIN1(n5918),
    .DIN1_t(n5918_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2047),
    .Q_t(WX2047_t)
  );


  nor2s3
  U3052
  (
    .DIN1(n5925),
    .DIN1_t(n5925_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2045),
    .Q_t(WX2045_t)
  );


  nor2s3
  U3053
  (
    .DIN1(n5932),
    .DIN1_t(n5932_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2043),
    .Q_t(WX2043_t)
  );


  nor2s3
  U3054
  (
    .DIN1(n5939),
    .DIN1_t(n5939_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2041),
    .Q_t(WX2041_t)
  );


  nor2s3
  U3055
  (
    .DIN1(n5946),
    .DIN1_t(n5946_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2039),
    .Q_t(WX2039_t)
  );


  nor2s3
  U3056
  (
    .DIN1(n5953),
    .DIN1_t(n5953_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2037),
    .Q_t(WX2037_t)
  );


  nor2s3
  U3057
  (
    .DIN1(n5960),
    .DIN1_t(n5960_t),
    .DIN2(n6759),
    .DIN2_t(n6759_t),
    .Q(WX2035),
    .Q_t(WX2035_t)
  );


  nor2s3
  U3058
  (
    .DIN1(n5967),
    .DIN1_t(n5967_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2033),
    .Q_t(WX2033_t)
  );


  nor2s3
  U3059
  (
    .DIN1(n5975),
    .DIN1_t(n5975_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2031),
    .Q_t(WX2031_t)
  );


  nor2s3
  U3060
  (
    .DIN1(n5984),
    .DIN1_t(n5984_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2029),
    .Q_t(WX2029_t)
  );


  nor2s3
  U3061
  (
    .DIN1(n5993),
    .DIN1_t(n5993_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2027),
    .Q_t(WX2027_t)
  );


  nor2s3
  U3062
  (
    .DIN1(n6002),
    .DIN1_t(n6002_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2025),
    .Q_t(WX2025_t)
  );


  nor2s3
  U3063
  (
    .DIN1(n6011),
    .DIN1_t(n6011_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2023),
    .Q_t(WX2023_t)
  );


  nor2s3
  U3064
  (
    .DIN1(n6020),
    .DIN1_t(n6020_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2021),
    .Q_t(WX2021_t)
  );


  nor2s3
  U3065
  (
    .DIN1(n6029),
    .DIN1_t(n6029_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2019),
    .Q_t(WX2019_t)
  );


  nor2s3
  U3066
  (
    .DIN1(n6038),
    .DIN1_t(n6038_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2017),
    .Q_t(WX2017_t)
  );


  nor2s3
  U3067
  (
    .DIN1(n6047),
    .DIN1_t(n6047_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2015),
    .Q_t(WX2015_t)
  );


  nor2s3
  U3068
  (
    .DIN1(n6056),
    .DIN1_t(n6056_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2013),
    .Q_t(WX2013_t)
  );


  nor2s3
  U3069
  (
    .DIN1(n6065),
    .DIN1_t(n6065_t),
    .DIN2(n6758),
    .DIN2_t(n6758_t),
    .Q(WX2011),
    .Q_t(WX2011_t)
  );


  nor2s3
  U3070
  (
    .DIN1(n6074),
    .DIN1_t(n6074_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX2009),
    .Q_t(WX2009_t)
  );


  nor2s3
  U3071
  (
    .DIN1(n6083),
    .DIN1_t(n6083_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX2007),
    .Q_t(WX2007_t)
  );


  nor2s3
  U3072
  (
    .DIN1(n6092),
    .DIN1_t(n6092_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX2005),
    .Q_t(WX2005_t)
  );


  nor2s3
  U3073
  (
    .DIN1(n6101),
    .DIN1_t(n6101_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX2003),
    .Q_t(WX2003_t)
  );


  nor2s3
  U3074
  (
    .DIN1(n6110),
    .DIN1_t(n6110_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX2001),
    .Q_t(WX2001_t)
  );


  nnd4s2
  U3075
  (
    .DIN1(n4234),
    .DIN1_t(n4234_t),
    .DIN2(n4235),
    .DIN2_t(n4235_t),
    .DIN3(n4236),
    .DIN3_t(n4236_t),
    .DIN4(n4237),
    .DIN4_t(n4237_t),
    .Q(WX1999),
    .Q_t(WX1999_t)
  );


  nnd2s3
  U3076
  (
    .DIN1(n3965),
    .DIN1_t(n3965_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4237),
    .Q_t(n4237_t)
  );


  xor2s3
  U3077
  (
    .DIN1(n4238),
    .DIN1_t(n4238_t),
    .DIN2(n4239),
    .DIN2_t(n4239_t),
    .Q(n3965),
    .Q_t(n3965_t)
  );


  xor2s3
  U3078
  (
    .DIN1(n5859),
    .DIN1_t(n5859_t),
    .DIN2(n5860),
    .DIN2_t(n5860_t),
    .Q(n4239),
    .Q_t(n4239_t)
  );


  xnr2s3
  U3079
  (
    .DIN1(n3285),
    .DIN1_t(n3285_t),
    .DIN2(n5861),
    .DIN2_t(n5861_t),
    .Q(n4238),
    .Q_t(n4238_t)
  );


  nnd2s3
  U3080
  (
    .DIN1(n3058),
    .DIN1_t(n3058_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4236),
    .Q_t(n4236_t)
  );


  xor2s3
  U3081
  (
    .DIN1(n4240),
    .DIN1_t(n4240_t),
    .DIN2(n4241),
    .DIN2_t(n4241_t),
    .Q(n3058),
    .Q_t(n3058_t)
  );


  xor2s3
  U3082
  (
    .DIN1(n5862),
    .DIN1_t(n5862_t),
    .DIN2(n5863),
    .DIN2_t(n5863_t),
    .Q(n4241),
    .Q_t(n4241_t)
  );


  xnr2s3
  U3083
  (
    .DIN1(n3286),
    .DIN1_t(n3286_t),
    .DIN2(n5864),
    .DIN2_t(n5864_t),
    .Q(n4240),
    .Q_t(n4240_t)
  );


  nnd2s3
  U3084
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2209),
    .DIN2_t(n2209_t),
    .Q(n4235),
    .Q_t(n4235_t)
  );


  nnd2s3
  U3085
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2208),
    .DIN2_t(n2208_t),
    .Q(n4234),
    .Q_t(n4234_t)
  );


  nnd4s2
  U3086
  (
    .DIN1(n4242),
    .DIN1_t(n4242_t),
    .DIN2(n4243),
    .DIN2_t(n4243_t),
    .DIN3(n4244),
    .DIN3_t(n4244_t),
    .DIN4(n4245),
    .DIN4_t(n4245_t),
    .Q(WX1997),
    .Q_t(WX1997_t)
  );


  nnd2s3
  U3087
  (
    .DIN1(n3972),
    .DIN1_t(n3972_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4245),
    .Q_t(n4245_t)
  );


  xor2s3
  U3088
  (
    .DIN1(n4246),
    .DIN1_t(n4246_t),
    .DIN2(n4247),
    .DIN2_t(n4247_t),
    .Q(n3972),
    .Q_t(n3972_t)
  );


  xor2s3
  U3089
  (
    .DIN1(n5866),
    .DIN1_t(n5866_t),
    .DIN2(n5867),
    .DIN2_t(n5867_t),
    .Q(n4247),
    .Q_t(n4247_t)
  );


  xnr2s3
  U3090
  (
    .DIN1(n3287),
    .DIN1_t(n3287_t),
    .DIN2(n5868),
    .DIN2_t(n5868_t),
    .Q(n4246),
    .Q_t(n4246_t)
  );


  nnd2s3
  U3091
  (
    .DIN1(n3064),
    .DIN1_t(n3064_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4244),
    .Q_t(n4244_t)
  );


  xor2s3
  U3092
  (
    .DIN1(n4248),
    .DIN1_t(n4248_t),
    .DIN2(n4249),
    .DIN2_t(n4249_t),
    .Q(n3064),
    .Q_t(n3064_t)
  );


  xor2s3
  U3093
  (
    .DIN1(n5869),
    .DIN1_t(n5869_t),
    .DIN2(n5870),
    .DIN2_t(n5870_t),
    .Q(n4249),
    .Q_t(n4249_t)
  );


  xnr2s3
  U3094
  (
    .DIN1(n3288),
    .DIN1_t(n3288_t),
    .DIN2(n5871),
    .DIN2_t(n5871_t),
    .Q(n4248),
    .Q_t(n4248_t)
  );


  nnd2s3
  U3095
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2210),
    .DIN2_t(n2210_t),
    .Q(n4243),
    .Q_t(n4243_t)
  );


  nnd2s3
  U3096
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2207),
    .DIN2_t(n2207_t),
    .Q(n4242),
    .Q_t(n4242_t)
  );


  nnd4s2
  U3097
  (
    .DIN1(n4250),
    .DIN1_t(n4250_t),
    .DIN2(n4251),
    .DIN2_t(n4251_t),
    .DIN3(n4252),
    .DIN3_t(n4252_t),
    .DIN4(n4253),
    .DIN4_t(n4253_t),
    .Q(WX1995),
    .Q_t(WX1995_t)
  );


  nnd2s3
  U3098
  (
    .DIN1(n3979),
    .DIN1_t(n3979_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4253),
    .Q_t(n4253_t)
  );


  xor2s3
  U3099
  (
    .DIN1(n4254),
    .DIN1_t(n4254_t),
    .DIN2(n4255),
    .DIN2_t(n4255_t),
    .Q(n3979),
    .Q_t(n3979_t)
  );


  xor2s3
  U3100
  (
    .DIN1(n5873),
    .DIN1_t(n5873_t),
    .DIN2(n5874),
    .DIN2_t(n5874_t),
    .Q(n4255),
    .Q_t(n4255_t)
  );


  xnr2s3
  U3101
  (
    .DIN1(n3289),
    .DIN1_t(n3289_t),
    .DIN2(n5875),
    .DIN2_t(n5875_t),
    .Q(n4254),
    .Q_t(n4254_t)
  );


  nnd2s3
  U3102
  (
    .DIN1(n3070),
    .DIN1_t(n3070_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4252),
    .Q_t(n4252_t)
  );


  xor2s3
  U3103
  (
    .DIN1(n4256),
    .DIN1_t(n4256_t),
    .DIN2(n4257),
    .DIN2_t(n4257_t),
    .Q(n3070),
    .Q_t(n3070_t)
  );


  xor2s3
  U3104
  (
    .DIN1(n5876),
    .DIN1_t(n5876_t),
    .DIN2(n5877),
    .DIN2_t(n5877_t),
    .Q(n4257),
    .Q_t(n4257_t)
  );


  xnr2s3
  U3105
  (
    .DIN1(n3290),
    .DIN1_t(n3290_t),
    .DIN2(n5878),
    .DIN2_t(n5878_t),
    .Q(n4256),
    .Q_t(n4256_t)
  );


  nnd2s3
  U3106
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2211),
    .DIN2_t(n2211_t),
    .Q(n4251),
    .Q_t(n4251_t)
  );


  nnd2s3
  U3107
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2206),
    .DIN2_t(n2206_t),
    .Q(n4250),
    .Q_t(n4250_t)
  );


  nnd4s2
  U3108
  (
    .DIN1(n4258),
    .DIN1_t(n4258_t),
    .DIN2(n4259),
    .DIN2_t(n4259_t),
    .DIN3(n4260),
    .DIN3_t(n4260_t),
    .DIN4(n4261),
    .DIN4_t(n4261_t),
    .Q(WX1993),
    .Q_t(WX1993_t)
  );


  nnd2s3
  U3109
  (
    .DIN1(n3986),
    .DIN1_t(n3986_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4261),
    .Q_t(n4261_t)
  );


  xor2s3
  U3110
  (
    .DIN1(n4262),
    .DIN1_t(n4262_t),
    .DIN2(n4263),
    .DIN2_t(n4263_t),
    .Q(n3986),
    .Q_t(n3986_t)
  );


  xor2s3
  U3111
  (
    .DIN1(n5880),
    .DIN1_t(n5880_t),
    .DIN2(n5881),
    .DIN2_t(n5881_t),
    .Q(n4263),
    .Q_t(n4263_t)
  );


  xnr2s3
  U3112
  (
    .DIN1(n3291),
    .DIN1_t(n3291_t),
    .DIN2(n5882),
    .DIN2_t(n5882_t),
    .Q(n4262),
    .Q_t(n4262_t)
  );


  nnd2s3
  U3113
  (
    .DIN1(n3076),
    .DIN1_t(n3076_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4260),
    .Q_t(n4260_t)
  );


  xor2s3
  U3114
  (
    .DIN1(n4264),
    .DIN1_t(n4264_t),
    .DIN2(n4265),
    .DIN2_t(n4265_t),
    .Q(n3076),
    .Q_t(n3076_t)
  );


  xor2s3
  U3115
  (
    .DIN1(n5883),
    .DIN1_t(n5883_t),
    .DIN2(n5884),
    .DIN2_t(n5884_t),
    .Q(n4265),
    .Q_t(n4265_t)
  );


  xnr2s3
  U3116
  (
    .DIN1(n3292),
    .DIN1_t(n3292_t),
    .DIN2(n5885),
    .DIN2_t(n5885_t),
    .Q(n4264),
    .Q_t(n4264_t)
  );


  nnd2s3
  U3117
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2212),
    .DIN2_t(n2212_t),
    .Q(n4259),
    .Q_t(n4259_t)
  );


  nnd2s3
  U3118
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2205),
    .DIN2_t(n2205_t),
    .Q(n4258),
    .Q_t(n4258_t)
  );


  nnd4s2
  U3119
  (
    .DIN1(n4266),
    .DIN1_t(n4266_t),
    .DIN2(n4267),
    .DIN2_t(n4267_t),
    .DIN3(n4268),
    .DIN3_t(n4268_t),
    .DIN4(n4269),
    .DIN4_t(n4269_t),
    .Q(WX1991),
    .Q_t(WX1991_t)
  );


  nnd2s3
  U3120
  (
    .DIN1(n3993),
    .DIN1_t(n3993_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4269),
    .Q_t(n4269_t)
  );


  xor2s3
  U3121
  (
    .DIN1(n4270),
    .DIN1_t(n4270_t),
    .DIN2(n4271),
    .DIN2_t(n4271_t),
    .Q(n3993),
    .Q_t(n3993_t)
  );


  xor2s3
  U3122
  (
    .DIN1(n5887),
    .DIN1_t(n5887_t),
    .DIN2(n5888),
    .DIN2_t(n5888_t),
    .Q(n4271),
    .Q_t(n4271_t)
  );


  xnr2s3
  U3123
  (
    .DIN1(n3293),
    .DIN1_t(n3293_t),
    .DIN2(n5889),
    .DIN2_t(n5889_t),
    .Q(n4270),
    .Q_t(n4270_t)
  );


  nnd2s3
  U3124
  (
    .DIN1(n3082),
    .DIN1_t(n3082_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4268),
    .Q_t(n4268_t)
  );


  xor2s3
  U3125
  (
    .DIN1(n4272),
    .DIN1_t(n4272_t),
    .DIN2(n4273),
    .DIN2_t(n4273_t),
    .Q(n3082),
    .Q_t(n3082_t)
  );


  xor2s3
  U3126
  (
    .DIN1(n5890),
    .DIN1_t(n5890_t),
    .DIN2(n5891),
    .DIN2_t(n5891_t),
    .Q(n4273),
    .Q_t(n4273_t)
  );


  xnr2s3
  U3127
  (
    .DIN1(n3294),
    .DIN1_t(n3294_t),
    .DIN2(n5892),
    .DIN2_t(n5892_t),
    .Q(n4272),
    .Q_t(n4272_t)
  );


  nnd2s3
  U3128
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2213),
    .DIN2_t(n2213_t),
    .Q(n4267),
    .Q_t(n4267_t)
  );


  nnd2s3
  U3129
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2204),
    .DIN2_t(n2204_t),
    .Q(n4266),
    .Q_t(n4266_t)
  );


  nnd4s2
  U3130
  (
    .DIN1(n4274),
    .DIN1_t(n4274_t),
    .DIN2(n4275),
    .DIN2_t(n4275_t),
    .DIN3(n4276),
    .DIN3_t(n4276_t),
    .DIN4(n4277),
    .DIN4_t(n4277_t),
    .Q(WX1989),
    .Q_t(WX1989_t)
  );


  nnd2s3
  U3131
  (
    .DIN1(n4000),
    .DIN1_t(n4000_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4277),
    .Q_t(n4277_t)
  );


  xor2s3
  U3132
  (
    .DIN1(n4278),
    .DIN1_t(n4278_t),
    .DIN2(n4279),
    .DIN2_t(n4279_t),
    .Q(n4000),
    .Q_t(n4000_t)
  );


  xor2s3
  U3133
  (
    .DIN1(n5894),
    .DIN1_t(n5894_t),
    .DIN2(n5895),
    .DIN2_t(n5895_t),
    .Q(n4279),
    .Q_t(n4279_t)
  );


  xnr2s3
  U3134
  (
    .DIN1(n3295),
    .DIN1_t(n3295_t),
    .DIN2(n5896),
    .DIN2_t(n5896_t),
    .Q(n4278),
    .Q_t(n4278_t)
  );


  nnd2s3
  U3135
  (
    .DIN1(n3088),
    .DIN1_t(n3088_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4276),
    .Q_t(n4276_t)
  );


  xor2s3
  U3136
  (
    .DIN1(n4280),
    .DIN1_t(n4280_t),
    .DIN2(n4281),
    .DIN2_t(n4281_t),
    .Q(n3088),
    .Q_t(n3088_t)
  );


  xor2s3
  U3137
  (
    .DIN1(n5897),
    .DIN1_t(n5897_t),
    .DIN2(n5898),
    .DIN2_t(n5898_t),
    .Q(n4281),
    .Q_t(n4281_t)
  );


  xnr2s3
  U3138
  (
    .DIN1(n3296),
    .DIN1_t(n3296_t),
    .DIN2(n5899),
    .DIN2_t(n5899_t),
    .Q(n4280),
    .Q_t(n4280_t)
  );


  nnd2s3
  U3139
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2214),
    .DIN2_t(n2214_t),
    .Q(n4275),
    .Q_t(n4275_t)
  );


  nnd2s3
  U3140
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2203),
    .DIN2_t(n2203_t),
    .Q(n4274),
    .Q_t(n4274_t)
  );


  nnd4s2
  U3141
  (
    .DIN1(n4282),
    .DIN1_t(n4282_t),
    .DIN2(n4283),
    .DIN2_t(n4283_t),
    .DIN3(n4284),
    .DIN3_t(n4284_t),
    .DIN4(n4285),
    .DIN4_t(n4285_t),
    .Q(WX1987),
    .Q_t(WX1987_t)
  );


  nnd2s3
  U3142
  (
    .DIN1(n4007),
    .DIN1_t(n4007_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4285),
    .Q_t(n4285_t)
  );


  xor2s3
  U3143
  (
    .DIN1(n4286),
    .DIN1_t(n4286_t),
    .DIN2(n4287),
    .DIN2_t(n4287_t),
    .Q(n4007),
    .Q_t(n4007_t)
  );


  xor2s3
  U3144
  (
    .DIN1(n5901),
    .DIN1_t(n5901_t),
    .DIN2(n5902),
    .DIN2_t(n5902_t),
    .Q(n4287),
    .Q_t(n4287_t)
  );


  xnr2s3
  U3145
  (
    .DIN1(n3297),
    .DIN1_t(n3297_t),
    .DIN2(n5903),
    .DIN2_t(n5903_t),
    .Q(n4286),
    .Q_t(n4286_t)
  );


  nnd2s3
  U3146
  (
    .DIN1(n3094),
    .DIN1_t(n3094_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4284),
    .Q_t(n4284_t)
  );


  xor2s3
  U3147
  (
    .DIN1(n4288),
    .DIN1_t(n4288_t),
    .DIN2(n4289),
    .DIN2_t(n4289_t),
    .Q(n3094),
    .Q_t(n3094_t)
  );


  xor2s3
  U3148
  (
    .DIN1(n5904),
    .DIN1_t(n5904_t),
    .DIN2(n5905),
    .DIN2_t(n5905_t),
    .Q(n4289),
    .Q_t(n4289_t)
  );


  xnr2s3
  U3149
  (
    .DIN1(n3298),
    .DIN1_t(n3298_t),
    .DIN2(n5906),
    .DIN2_t(n5906_t),
    .Q(n4288),
    .Q_t(n4288_t)
  );


  nnd2s3
  U3150
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2215),
    .DIN2_t(n2215_t),
    .Q(n4283),
    .Q_t(n4283_t)
  );


  nnd2s3
  U3151
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2202),
    .DIN2_t(n2202_t),
    .Q(n4282),
    .Q_t(n4282_t)
  );


  nnd4s2
  U3152
  (
    .DIN1(n4290),
    .DIN1_t(n4290_t),
    .DIN2(n4291),
    .DIN2_t(n4291_t),
    .DIN3(n4292),
    .DIN3_t(n4292_t),
    .DIN4(n4293),
    .DIN4_t(n4293_t),
    .Q(WX1985),
    .Q_t(WX1985_t)
  );


  nnd2s3
  U3153
  (
    .DIN1(n4014),
    .DIN1_t(n4014_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4293),
    .Q_t(n4293_t)
  );


  xor2s3
  U3154
  (
    .DIN1(n4294),
    .DIN1_t(n4294_t),
    .DIN2(n4295),
    .DIN2_t(n4295_t),
    .Q(n4014),
    .Q_t(n4014_t)
  );


  xor2s3
  U3155
  (
    .DIN1(n5908),
    .DIN1_t(n5908_t),
    .DIN2(n5909),
    .DIN2_t(n5909_t),
    .Q(n4295),
    .Q_t(n4295_t)
  );


  xnr2s3
  U3156
  (
    .DIN1(n3299),
    .DIN1_t(n3299_t),
    .DIN2(n5910),
    .DIN2_t(n5910_t),
    .Q(n4294),
    .Q_t(n4294_t)
  );


  nnd2s3
  U3157
  (
    .DIN1(n3100),
    .DIN1_t(n3100_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4292),
    .Q_t(n4292_t)
  );


  xor2s3
  U3158
  (
    .DIN1(n4296),
    .DIN1_t(n4296_t),
    .DIN2(n4297),
    .DIN2_t(n4297_t),
    .Q(n3100),
    .Q_t(n3100_t)
  );


  xor2s3
  U3159
  (
    .DIN1(n5911),
    .DIN1_t(n5911_t),
    .DIN2(n5912),
    .DIN2_t(n5912_t),
    .Q(n4297),
    .Q_t(n4297_t)
  );


  xnr2s3
  U3160
  (
    .DIN1(n3300),
    .DIN1_t(n3300_t),
    .DIN2(n5913),
    .DIN2_t(n5913_t),
    .Q(n4296),
    .Q_t(n4296_t)
  );


  nnd2s3
  U3161
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2216),
    .DIN2_t(n2216_t),
    .Q(n4291),
    .Q_t(n4291_t)
  );


  nnd2s3
  U3162
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2201),
    .DIN2_t(n2201_t),
    .Q(n4290),
    .Q_t(n4290_t)
  );


  nnd4s2
  U3163
  (
    .DIN1(n4298),
    .DIN1_t(n4298_t),
    .DIN2(n4299),
    .DIN2_t(n4299_t),
    .DIN3(n4300),
    .DIN3_t(n4300_t),
    .DIN4(n4301),
    .DIN4_t(n4301_t),
    .Q(WX1983),
    .Q_t(WX1983_t)
  );


  nnd2s3
  U3164
  (
    .DIN1(n4021),
    .DIN1_t(n4021_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4301),
    .Q_t(n4301_t)
  );


  xor2s3
  U3165
  (
    .DIN1(n4302),
    .DIN1_t(n4302_t),
    .DIN2(n4303),
    .DIN2_t(n4303_t),
    .Q(n4021),
    .Q_t(n4021_t)
  );


  xor2s3
  U3166
  (
    .DIN1(n5915),
    .DIN1_t(n5915_t),
    .DIN2(n5916),
    .DIN2_t(n5916_t),
    .Q(n4303),
    .Q_t(n4303_t)
  );


  xnr2s3
  U3167
  (
    .DIN1(n3301),
    .DIN1_t(n3301_t),
    .DIN2(n5917),
    .DIN2_t(n5917_t),
    .Q(n4302),
    .Q_t(n4302_t)
  );


  nnd2s3
  U3168
  (
    .DIN1(n3106),
    .DIN1_t(n3106_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4300),
    .Q_t(n4300_t)
  );


  xor2s3
  U3169
  (
    .DIN1(n4304),
    .DIN1_t(n4304_t),
    .DIN2(n4305),
    .DIN2_t(n4305_t),
    .Q(n3106),
    .Q_t(n3106_t)
  );


  xor2s3
  U3170
  (
    .DIN1(n5918),
    .DIN1_t(n5918_t),
    .DIN2(n5919),
    .DIN2_t(n5919_t),
    .Q(n4305),
    .Q_t(n4305_t)
  );


  xnr2s3
  U3171
  (
    .DIN1(n3302),
    .DIN1_t(n3302_t),
    .DIN2(n5920),
    .DIN2_t(n5920_t),
    .Q(n4304),
    .Q_t(n4304_t)
  );


  nnd2s3
  U3172
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2217),
    .DIN2_t(n2217_t),
    .Q(n4299),
    .Q_t(n4299_t)
  );


  nnd2s3
  U3173
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2200),
    .DIN2_t(n2200_t),
    .Q(n4298),
    .Q_t(n4298_t)
  );


  nnd4s2
  U3174
  (
    .DIN1(n4306),
    .DIN1_t(n4306_t),
    .DIN2(n4307),
    .DIN2_t(n4307_t),
    .DIN3(n4308),
    .DIN3_t(n4308_t),
    .DIN4(n4309),
    .DIN4_t(n4309_t),
    .Q(WX1981),
    .Q_t(WX1981_t)
  );


  nnd2s3
  U3175
  (
    .DIN1(n4028),
    .DIN1_t(n4028_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4309),
    .Q_t(n4309_t)
  );


  xor2s3
  U3176
  (
    .DIN1(n4310),
    .DIN1_t(n4310_t),
    .DIN2(n4311),
    .DIN2_t(n4311_t),
    .Q(n4028),
    .Q_t(n4028_t)
  );


  xor2s3
  U3177
  (
    .DIN1(n5922),
    .DIN1_t(n5922_t),
    .DIN2(n5923),
    .DIN2_t(n5923_t),
    .Q(n4311),
    .Q_t(n4311_t)
  );


  xnr2s3
  U3178
  (
    .DIN1(n3303),
    .DIN1_t(n3303_t),
    .DIN2(n5924),
    .DIN2_t(n5924_t),
    .Q(n4310),
    .Q_t(n4310_t)
  );


  nnd2s3
  U3179
  (
    .DIN1(n3112),
    .DIN1_t(n3112_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4308),
    .Q_t(n4308_t)
  );


  xor2s3
  U3180
  (
    .DIN1(n4312),
    .DIN1_t(n4312_t),
    .DIN2(n4313),
    .DIN2_t(n4313_t),
    .Q(n3112),
    .Q_t(n3112_t)
  );


  xor2s3
  U3181
  (
    .DIN1(n5925),
    .DIN1_t(n5925_t),
    .DIN2(n5926),
    .DIN2_t(n5926_t),
    .Q(n4313),
    .Q_t(n4313_t)
  );


  xnr2s3
  U3182
  (
    .DIN1(n3304),
    .DIN1_t(n3304_t),
    .DIN2(n5927),
    .DIN2_t(n5927_t),
    .Q(n4312),
    .Q_t(n4312_t)
  );


  nnd2s3
  U3183
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2218),
    .DIN2_t(n2218_t),
    .Q(n4307),
    .Q_t(n4307_t)
  );


  nnd2s3
  U3184
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2199),
    .DIN2_t(n2199_t),
    .Q(n4306),
    .Q_t(n4306_t)
  );


  nnd4s2
  U3185
  (
    .DIN1(n4314),
    .DIN1_t(n4314_t),
    .DIN2(n4315),
    .DIN2_t(n4315_t),
    .DIN3(n4316),
    .DIN3_t(n4316_t),
    .DIN4(n4317),
    .DIN4_t(n4317_t),
    .Q(WX1979),
    .Q_t(WX1979_t)
  );


  nnd2s3
  U3186
  (
    .DIN1(n4035),
    .DIN1_t(n4035_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4317),
    .Q_t(n4317_t)
  );


  xor2s3
  U3187
  (
    .DIN1(n4318),
    .DIN1_t(n4318_t),
    .DIN2(n4319),
    .DIN2_t(n4319_t),
    .Q(n4035),
    .Q_t(n4035_t)
  );


  xor2s3
  U3188
  (
    .DIN1(n5929),
    .DIN1_t(n5929_t),
    .DIN2(n5930),
    .DIN2_t(n5930_t),
    .Q(n4319),
    .Q_t(n4319_t)
  );


  xnr2s3
  U3189
  (
    .DIN1(n3305),
    .DIN1_t(n3305_t),
    .DIN2(n5931),
    .DIN2_t(n5931_t),
    .Q(n4318),
    .Q_t(n4318_t)
  );


  nnd2s3
  U3190
  (
    .DIN1(n3118),
    .DIN1_t(n3118_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4316),
    .Q_t(n4316_t)
  );


  xor2s3
  U3191
  (
    .DIN1(n4320),
    .DIN1_t(n4320_t),
    .DIN2(n4321),
    .DIN2_t(n4321_t),
    .Q(n3118),
    .Q_t(n3118_t)
  );


  xor2s3
  U3192
  (
    .DIN1(n5932),
    .DIN1_t(n5932_t),
    .DIN2(n5933),
    .DIN2_t(n5933_t),
    .Q(n4321),
    .Q_t(n4321_t)
  );


  xnr2s3
  U3193
  (
    .DIN1(n3306),
    .DIN1_t(n3306_t),
    .DIN2(n5934),
    .DIN2_t(n5934_t),
    .Q(n4320),
    .Q_t(n4320_t)
  );


  nnd2s3
  U3194
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2219),
    .DIN2_t(n2219_t),
    .Q(n4315),
    .Q_t(n4315_t)
  );


  nnd2s3
  U3195
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2198),
    .DIN2_t(n2198_t),
    .Q(n4314),
    .Q_t(n4314_t)
  );


  nnd4s2
  U3196
  (
    .DIN1(n4322),
    .DIN1_t(n4322_t),
    .DIN2(n4323),
    .DIN2_t(n4323_t),
    .DIN3(n4324),
    .DIN3_t(n4324_t),
    .DIN4(n4325),
    .DIN4_t(n4325_t),
    .Q(WX1977),
    .Q_t(WX1977_t)
  );


  nnd2s3
  U3197
  (
    .DIN1(n4042),
    .DIN1_t(n4042_t),
    .DIN2(n6640),
    .DIN2_t(n6640_t),
    .Q(n4325),
    .Q_t(n4325_t)
  );


  xor2s3
  U3198
  (
    .DIN1(n4326),
    .DIN1_t(n4326_t),
    .DIN2(n4327),
    .DIN2_t(n4327_t),
    .Q(n4042),
    .Q_t(n4042_t)
  );


  xor2s3
  U3199
  (
    .DIN1(n5936),
    .DIN1_t(n5936_t),
    .DIN2(n5937),
    .DIN2_t(n5937_t),
    .Q(n4327),
    .Q_t(n4327_t)
  );


  xnr2s3
  U3200
  (
    .DIN1(n3307),
    .DIN1_t(n3307_t),
    .DIN2(n5938),
    .DIN2_t(n5938_t),
    .Q(n4326),
    .Q_t(n4326_t)
  );


  nnd2s3
  U3201
  (
    .DIN1(n3124),
    .DIN1_t(n3124_t),
    .DIN2(n6671),
    .DIN2_t(n6671_t),
    .Q(n4324),
    .Q_t(n4324_t)
  );


  xor2s3
  U3202
  (
    .DIN1(n4328),
    .DIN1_t(n4328_t),
    .DIN2(n4329),
    .DIN2_t(n4329_t),
    .Q(n3124),
    .Q_t(n3124_t)
  );


  xor2s3
  U3203
  (
    .DIN1(n5939),
    .DIN1_t(n5939_t),
    .DIN2(n5940),
    .DIN2_t(n5940_t),
    .Q(n4329),
    .Q_t(n4329_t)
  );


  xnr2s3
  U3204
  (
    .DIN1(n3308),
    .DIN1_t(n3308_t),
    .DIN2(n5941),
    .DIN2_t(n5941_t),
    .Q(n4328),
    .Q_t(n4328_t)
  );


  nnd2s3
  U3205
  (
    .DIN1(n6598),
    .DIN1_t(n6598_t),
    .DIN2(n2220),
    .DIN2_t(n2220_t),
    .Q(n4323),
    .Q_t(n4323_t)
  );


  nnd2s3
  U3206
  (
    .DIN1(n6567),
    .DIN1_t(n6567_t),
    .DIN2(n2197),
    .DIN2_t(n2197_t),
    .Q(n4322),
    .Q_t(n4322_t)
  );


  nnd4s2
  U3207
  (
    .DIN1(n4330),
    .DIN1_t(n4330_t),
    .DIN2(n4331),
    .DIN2_t(n4331_t),
    .DIN3(n4332),
    .DIN3_t(n4332_t),
    .DIN4(n4333),
    .DIN4_t(n4333_t),
    .Q(WX1975),
    .Q_t(WX1975_t)
  );


  nnd2s3
  U3208
  (
    .DIN1(n4049),
    .DIN1_t(n4049_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4333),
    .Q_t(n4333_t)
  );


  xor2s3
  U3209
  (
    .DIN1(n4334),
    .DIN1_t(n4334_t),
    .DIN2(n4335),
    .DIN2_t(n4335_t),
    .Q(n4049),
    .Q_t(n4049_t)
  );


  xor2s3
  U3210
  (
    .DIN1(n5943),
    .DIN1_t(n5943_t),
    .DIN2(n5944),
    .DIN2_t(n5944_t),
    .Q(n4335),
    .Q_t(n4335_t)
  );


  xnr2s3
  U3211
  (
    .DIN1(n3309),
    .DIN1_t(n3309_t),
    .DIN2(n5945),
    .DIN2_t(n5945_t),
    .Q(n4334),
    .Q_t(n4334_t)
  );


  nnd2s3
  U3212
  (
    .DIN1(n3130),
    .DIN1_t(n3130_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4332),
    .Q_t(n4332_t)
  );


  xor2s3
  U3213
  (
    .DIN1(n4336),
    .DIN1_t(n4336_t),
    .DIN2(n4337),
    .DIN2_t(n4337_t),
    .Q(n3130),
    .Q_t(n3130_t)
  );


  xor2s3
  U3214
  (
    .DIN1(n5946),
    .DIN1_t(n5946_t),
    .DIN2(n5947),
    .DIN2_t(n5947_t),
    .Q(n4337),
    .Q_t(n4337_t)
  );


  xnr2s3
  U3215
  (
    .DIN1(n3310),
    .DIN1_t(n3310_t),
    .DIN2(n5948),
    .DIN2_t(n5948_t),
    .Q(n4336),
    .Q_t(n4336_t)
  );


  nnd2s3
  U3216
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2221),
    .DIN2_t(n2221_t),
    .Q(n4331),
    .Q_t(n4331_t)
  );


  nnd2s3
  U3217
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2196),
    .DIN2_t(n2196_t),
    .Q(n4330),
    .Q_t(n4330_t)
  );


  nnd4s2
  U3218
  (
    .DIN1(n4338),
    .DIN1_t(n4338_t),
    .DIN2(n4339),
    .DIN2_t(n4339_t),
    .DIN3(n4340),
    .DIN3_t(n4340_t),
    .DIN4(n4341),
    .DIN4_t(n4341_t),
    .Q(WX1973),
    .Q_t(WX1973_t)
  );


  nnd2s3
  U3219
  (
    .DIN1(n4056),
    .DIN1_t(n4056_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4341),
    .Q_t(n4341_t)
  );


  xor2s3
  U3220
  (
    .DIN1(n4342),
    .DIN1_t(n4342_t),
    .DIN2(n4343),
    .DIN2_t(n4343_t),
    .Q(n4056),
    .Q_t(n4056_t)
  );


  xor2s3
  U3221
  (
    .DIN1(n5950),
    .DIN1_t(n5950_t),
    .DIN2(n5951),
    .DIN2_t(n5951_t),
    .Q(n4343),
    .Q_t(n4343_t)
  );


  xnr2s3
  U3222
  (
    .DIN1(n3311),
    .DIN1_t(n3311_t),
    .DIN2(n5952),
    .DIN2_t(n5952_t),
    .Q(n4342),
    .Q_t(n4342_t)
  );


  nnd2s3
  U3223
  (
    .DIN1(n3136),
    .DIN1_t(n3136_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4340),
    .Q_t(n4340_t)
  );


  xor2s3
  U3224
  (
    .DIN1(n4344),
    .DIN1_t(n4344_t),
    .DIN2(n4345),
    .DIN2_t(n4345_t),
    .Q(n3136),
    .Q_t(n3136_t)
  );


  xor2s3
  U3225
  (
    .DIN1(n5953),
    .DIN1_t(n5953_t),
    .DIN2(n5954),
    .DIN2_t(n5954_t),
    .Q(n4345),
    .Q_t(n4345_t)
  );


  xnr2s3
  U3226
  (
    .DIN1(n3312),
    .DIN1_t(n3312_t),
    .DIN2(n5955),
    .DIN2_t(n5955_t),
    .Q(n4344),
    .Q_t(n4344_t)
  );


  nnd2s3
  U3227
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2222),
    .DIN2_t(n2222_t),
    .Q(n4339),
    .Q_t(n4339_t)
  );


  nnd2s3
  U3228
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2195),
    .DIN2_t(n2195_t),
    .Q(n4338),
    .Q_t(n4338_t)
  );


  nnd4s2
  U3229
  (
    .DIN1(n4346),
    .DIN1_t(n4346_t),
    .DIN2(n4347),
    .DIN2_t(n4347_t),
    .DIN3(n4348),
    .DIN3_t(n4348_t),
    .DIN4(n4349),
    .DIN4_t(n4349_t),
    .Q(WX1971),
    .Q_t(WX1971_t)
  );


  nnd2s3
  U3230
  (
    .DIN1(n4063),
    .DIN1_t(n4063_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4349),
    .Q_t(n4349_t)
  );


  xor2s3
  U3231
  (
    .DIN1(n4350),
    .DIN1_t(n4350_t),
    .DIN2(n4351),
    .DIN2_t(n4351_t),
    .Q(n4063),
    .Q_t(n4063_t)
  );


  xor2s3
  U3232
  (
    .DIN1(n5957),
    .DIN1_t(n5957_t),
    .DIN2(n5958),
    .DIN2_t(n5958_t),
    .Q(n4351),
    .Q_t(n4351_t)
  );


  xnr2s3
  U3233
  (
    .DIN1(n3313),
    .DIN1_t(n3313_t),
    .DIN2(n5959),
    .DIN2_t(n5959_t),
    .Q(n4350),
    .Q_t(n4350_t)
  );


  nnd2s3
  U3234
  (
    .DIN1(n3142),
    .DIN1_t(n3142_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4348),
    .Q_t(n4348_t)
  );


  xor2s3
  U3235
  (
    .DIN1(n4352),
    .DIN1_t(n4352_t),
    .DIN2(n4353),
    .DIN2_t(n4353_t),
    .Q(n3142),
    .Q_t(n3142_t)
  );


  xor2s3
  U3236
  (
    .DIN1(n5960),
    .DIN1_t(n5960_t),
    .DIN2(n5961),
    .DIN2_t(n5961_t),
    .Q(n4353),
    .Q_t(n4353_t)
  );


  xnr2s3
  U3237
  (
    .DIN1(n3314),
    .DIN1_t(n3314_t),
    .DIN2(n5962),
    .DIN2_t(n5962_t),
    .Q(n4352),
    .Q_t(n4352_t)
  );


  nnd2s3
  U3238
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2223),
    .DIN2_t(n2223_t),
    .Q(n4347),
    .Q_t(n4347_t)
  );


  nnd2s3
  U3239
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2194),
    .DIN2_t(n2194_t),
    .Q(n4346),
    .Q_t(n4346_t)
  );


  nnd4s2
  U3240
  (
    .DIN1(n4354),
    .DIN1_t(n4354_t),
    .DIN2(n4355),
    .DIN2_t(n4355_t),
    .DIN3(n4356),
    .DIN3_t(n4356_t),
    .DIN4(n4357),
    .DIN4_t(n4357_t),
    .Q(WX1969),
    .Q_t(WX1969_t)
  );


  nnd2s3
  U3241
  (
    .DIN1(n4070),
    .DIN1_t(n4070_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4357),
    .Q_t(n4357_t)
  );


  xor2s3
  U3242
  (
    .DIN1(n4358),
    .DIN1_t(n4358_t),
    .DIN2(n4359),
    .DIN2_t(n4359_t),
    .Q(n4070),
    .Q_t(n4070_t)
  );


  xor2s3
  U3243
  (
    .DIN1(n5964),
    .DIN1_t(n5964_t),
    .DIN2(n5965),
    .DIN2_t(n5965_t),
    .Q(n4359),
    .Q_t(n4359_t)
  );


  xnr2s3
  U3244
  (
    .DIN1(n3315),
    .DIN1_t(n3315_t),
    .DIN2(n5966),
    .DIN2_t(n5966_t),
    .Q(n4358),
    .Q_t(n4358_t)
  );


  nnd2s3
  U3245
  (
    .DIN1(n3148),
    .DIN1_t(n3148_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4356),
    .Q_t(n4356_t)
  );


  xor2s3
  U3246
  (
    .DIN1(n4360),
    .DIN1_t(n4360_t),
    .DIN2(n4361),
    .DIN2_t(n4361_t),
    .Q(n3148),
    .Q_t(n3148_t)
  );


  xor2s3
  U3247
  (
    .DIN1(n5967),
    .DIN1_t(n5967_t),
    .DIN2(n5968),
    .DIN2_t(n5968_t),
    .Q(n4361),
    .Q_t(n4361_t)
  );


  xnr2s3
  U3248
  (
    .DIN1(n3316),
    .DIN1_t(n3316_t),
    .DIN2(n5969),
    .DIN2_t(n5969_t),
    .Q(n4360),
    .Q_t(n4360_t)
  );


  nnd2s3
  U3249
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2224),
    .DIN2_t(n2224_t),
    .Q(n4355),
    .Q_t(n4355_t)
  );


  nnd2s3
  U3250
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2193),
    .DIN2_t(n2193_t),
    .Q(n4354),
    .Q_t(n4354_t)
  );


  nnd4s2
  U3251
  (
    .DIN1(n4362),
    .DIN1_t(n4362_t),
    .DIN2(n4363),
    .DIN2_t(n4363_t),
    .DIN3(n4364),
    .DIN3_t(n4364_t),
    .DIN4(n4365),
    .DIN4_t(n4365_t),
    .Q(WX1967),
    .Q_t(WX1967_t)
  );


  nnd2s3
  U3252
  (
    .DIN1(n4078),
    .DIN1_t(n4078_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4365),
    .Q_t(n4365_t)
  );


  xor2s3
  U3253
  (
    .DIN1(n4366),
    .DIN1_t(n4366_t),
    .DIN2(n4367),
    .DIN2_t(n4367_t),
    .Q(n4078),
    .Q_t(n4078_t)
  );


  xor2s3
  U3254
  (
    .DIN1(n5973),
    .DIN1_t(n5973_t),
    .DIN2(n4368),
    .DIN2_t(n4368_t),
    .Q(n4367),
    .Q_t(n4367_t)
  );


  xor2s3
  U3255
  (
    .DIN1(n5971),
    .DIN1_t(n5971_t),
    .DIN2(n5972),
    .DIN2_t(n5972_t),
    .Q(n4368),
    .Q_t(n4368_t)
  );


  xor2s3
  U3256
  (
    .DIN1(n5974),
    .DIN1_t(n5974_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4366),
    .Q_t(n4366_t)
  );


  nnd2s3
  U3257
  (
    .DIN1(n3154),
    .DIN1_t(n3154_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4364),
    .Q_t(n4364_t)
  );


  xor2s3
  U3258
  (
    .DIN1(n4369),
    .DIN1_t(n4369_t),
    .DIN2(n4370),
    .DIN2_t(n4370_t),
    .Q(n3154),
    .Q_t(n3154_t)
  );


  xor2s3
  U3259
  (
    .DIN1(n5977),
    .DIN1_t(n5977_t),
    .DIN2(n4371),
    .DIN2_t(n4371_t),
    .Q(n4370),
    .Q_t(n4370_t)
  );


  xor2s3
  U3260
  (
    .DIN1(n5975),
    .DIN1_t(n5975_t),
    .DIN2(n5976),
    .DIN2_t(n5976_t),
    .Q(n4371),
    .Q_t(n4371_t)
  );


  xor2s3
  U3261
  (
    .DIN1(n5978),
    .DIN1_t(n5978_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4369),
    .Q_t(n4369_t)
  );


  nnd2s3
  U3262
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2225),
    .DIN2_t(n2225_t),
    .Q(n4363),
    .Q_t(n4363_t)
  );


  nnd2s3
  U3263
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2192),
    .DIN2_t(n2192_t),
    .Q(n4362),
    .Q_t(n4362_t)
  );


  nnd4s2
  U3264
  (
    .DIN1(n4372),
    .DIN1_t(n4372_t),
    .DIN2(n4373),
    .DIN2_t(n4373_t),
    .DIN3(n4374),
    .DIN3_t(n4374_t),
    .DIN4(n4375),
    .DIN4_t(n4375_t),
    .Q(WX1965),
    .Q_t(WX1965_t)
  );


  nnd2s3
  U3265
  (
    .DIN1(n4086),
    .DIN1_t(n4086_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4375),
    .Q_t(n4375_t)
  );


  xor2s3
  U3266
  (
    .DIN1(n4376),
    .DIN1_t(n4376_t),
    .DIN2(n4377),
    .DIN2_t(n4377_t),
    .Q(n4086),
    .Q_t(n4086_t)
  );


  xor2s3
  U3267
  (
    .DIN1(n5982),
    .DIN1_t(n5982_t),
    .DIN2(n4378),
    .DIN2_t(n4378_t),
    .Q(n4377),
    .Q_t(n4377_t)
  );


  xor2s3
  U3268
  (
    .DIN1(n5980),
    .DIN1_t(n5980_t),
    .DIN2(n5981),
    .DIN2_t(n5981_t),
    .Q(n4378),
    .Q_t(n4378_t)
  );


  xor2s3
  U3269
  (
    .DIN1(n5983),
    .DIN1_t(n5983_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4376),
    .Q_t(n4376_t)
  );


  nnd2s3
  U3270
  (
    .DIN1(n3160),
    .DIN1_t(n3160_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4374),
    .Q_t(n4374_t)
  );


  xor2s3
  U3271
  (
    .DIN1(n4379),
    .DIN1_t(n4379_t),
    .DIN2(n4380),
    .DIN2_t(n4380_t),
    .Q(n3160),
    .Q_t(n3160_t)
  );


  xor2s3
  U3272
  (
    .DIN1(n5986),
    .DIN1_t(n5986_t),
    .DIN2(n4381),
    .DIN2_t(n4381_t),
    .Q(n4380),
    .Q_t(n4380_t)
  );


  xor2s3
  U3273
  (
    .DIN1(n5984),
    .DIN1_t(n5984_t),
    .DIN2(n5985),
    .DIN2_t(n5985_t),
    .Q(n4381),
    .Q_t(n4381_t)
  );


  xor2s3
  U3274
  (
    .DIN1(n5987),
    .DIN1_t(n5987_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4379),
    .Q_t(n4379_t)
  );


  nnd2s3
  U3275
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2226),
    .DIN2_t(n2226_t),
    .Q(n4373),
    .Q_t(n4373_t)
  );


  nnd2s3
  U3276
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2191),
    .DIN2_t(n2191_t),
    .Q(n4372),
    .Q_t(n4372_t)
  );


  nnd4s2
  U3277
  (
    .DIN1(n4382),
    .DIN1_t(n4382_t),
    .DIN2(n4383),
    .DIN2_t(n4383_t),
    .DIN3(n4384),
    .DIN3_t(n4384_t),
    .DIN4(n4385),
    .DIN4_t(n4385_t),
    .Q(WX1963),
    .Q_t(WX1963_t)
  );


  nnd2s3
  U3278
  (
    .DIN1(n4094),
    .DIN1_t(n4094_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4385),
    .Q_t(n4385_t)
  );


  xor2s3
  U3279
  (
    .DIN1(n4386),
    .DIN1_t(n4386_t),
    .DIN2(n4387),
    .DIN2_t(n4387_t),
    .Q(n4094),
    .Q_t(n4094_t)
  );


  xor2s3
  U3280
  (
    .DIN1(n5991),
    .DIN1_t(n5991_t),
    .DIN2(n4388),
    .DIN2_t(n4388_t),
    .Q(n4387),
    .Q_t(n4387_t)
  );


  xor2s3
  U3281
  (
    .DIN1(n5989),
    .DIN1_t(n5989_t),
    .DIN2(n5990),
    .DIN2_t(n5990_t),
    .Q(n4388),
    .Q_t(n4388_t)
  );


  xor2s3
  U3282
  (
    .DIN1(n5992),
    .DIN1_t(n5992_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4386),
    .Q_t(n4386_t)
  );


  nnd2s3
  U3283
  (
    .DIN1(n3166),
    .DIN1_t(n3166_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4384),
    .Q_t(n4384_t)
  );


  xor2s3
  U3284
  (
    .DIN1(n4389),
    .DIN1_t(n4389_t),
    .DIN2(n4390),
    .DIN2_t(n4390_t),
    .Q(n3166),
    .Q_t(n3166_t)
  );


  xor2s3
  U3285
  (
    .DIN1(n5995),
    .DIN1_t(n5995_t),
    .DIN2(n4391),
    .DIN2_t(n4391_t),
    .Q(n4390),
    .Q_t(n4390_t)
  );


  xor2s3
  U3286
  (
    .DIN1(n5993),
    .DIN1_t(n5993_t),
    .DIN2(n5994),
    .DIN2_t(n5994_t),
    .Q(n4391),
    .Q_t(n4391_t)
  );


  xor2s3
  U3287
  (
    .DIN1(n5996),
    .DIN1_t(n5996_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4389),
    .Q_t(n4389_t)
  );


  nnd2s3
  U3288
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2227),
    .DIN2_t(n2227_t),
    .Q(n4383),
    .Q_t(n4383_t)
  );


  nnd2s3
  U3289
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2190),
    .DIN2_t(n2190_t),
    .Q(n4382),
    .Q_t(n4382_t)
  );


  nnd4s2
  U3290
  (
    .DIN1(n4392),
    .DIN1_t(n4392_t),
    .DIN2(n4393),
    .DIN2_t(n4393_t),
    .DIN3(n4394),
    .DIN3_t(n4394_t),
    .DIN4(n4395),
    .DIN4_t(n4395_t),
    .Q(WX1961),
    .Q_t(WX1961_t)
  );


  nnd2s3
  U3291
  (
    .DIN1(n4102),
    .DIN1_t(n4102_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4395),
    .Q_t(n4395_t)
  );


  xor2s3
  U3292
  (
    .DIN1(n4396),
    .DIN1_t(n4396_t),
    .DIN2(n4397),
    .DIN2_t(n4397_t),
    .Q(n4102),
    .Q_t(n4102_t)
  );


  xor2s3
  U3293
  (
    .DIN1(n6000),
    .DIN1_t(n6000_t),
    .DIN2(n4398),
    .DIN2_t(n4398_t),
    .Q(n4397),
    .Q_t(n4397_t)
  );


  xor2s3
  U3294
  (
    .DIN1(n5998),
    .DIN1_t(n5998_t),
    .DIN2(n5999),
    .DIN2_t(n5999_t),
    .Q(n4398),
    .Q_t(n4398_t)
  );


  xor2s3
  U3295
  (
    .DIN1(n6001),
    .DIN1_t(n6001_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4396),
    .Q_t(n4396_t)
  );


  nnd2s3
  U3296
  (
    .DIN1(n3172),
    .DIN1_t(n3172_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4394),
    .Q_t(n4394_t)
  );


  xor2s3
  U3297
  (
    .DIN1(n4399),
    .DIN1_t(n4399_t),
    .DIN2(n4400),
    .DIN2_t(n4400_t),
    .Q(n3172),
    .Q_t(n3172_t)
  );


  xor2s3
  U3298
  (
    .DIN1(n6004),
    .DIN1_t(n6004_t),
    .DIN2(n4401),
    .DIN2_t(n4401_t),
    .Q(n4400),
    .Q_t(n4400_t)
  );


  xor2s3
  U3299
  (
    .DIN1(n6002),
    .DIN1_t(n6002_t),
    .DIN2(n6003),
    .DIN2_t(n6003_t),
    .Q(n4401),
    .Q_t(n4401_t)
  );


  xor2s3
  U3300
  (
    .DIN1(n6005),
    .DIN1_t(n6005_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4399),
    .Q_t(n4399_t)
  );


  nnd2s3
  U3301
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2228),
    .DIN2_t(n2228_t),
    .Q(n4393),
    .Q_t(n4393_t)
  );


  nnd2s3
  U3302
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2189),
    .DIN2_t(n2189_t),
    .Q(n4392),
    .Q_t(n4392_t)
  );


  nnd4s2
  U3303
  (
    .DIN1(n4402),
    .DIN1_t(n4402_t),
    .DIN2(n4403),
    .DIN2_t(n4403_t),
    .DIN3(n4404),
    .DIN3_t(n4404_t),
    .DIN4(n4405),
    .DIN4_t(n4405_t),
    .Q(WX1959),
    .Q_t(WX1959_t)
  );


  nnd2s3
  U3304
  (
    .DIN1(n4110),
    .DIN1_t(n4110_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4405),
    .Q_t(n4405_t)
  );


  xor2s3
  U3305
  (
    .DIN1(n4406),
    .DIN1_t(n4406_t),
    .DIN2(n4407),
    .DIN2_t(n4407_t),
    .Q(n4110),
    .Q_t(n4110_t)
  );


  xor2s3
  U3306
  (
    .DIN1(n6009),
    .DIN1_t(n6009_t),
    .DIN2(n4408),
    .DIN2_t(n4408_t),
    .Q(n4407),
    .Q_t(n4407_t)
  );


  xor2s3
  U3307
  (
    .DIN1(n6007),
    .DIN1_t(n6007_t),
    .DIN2(n6008),
    .DIN2_t(n6008_t),
    .Q(n4408),
    .Q_t(n4408_t)
  );


  xor2s3
  U3308
  (
    .DIN1(n6010),
    .DIN1_t(n6010_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4406),
    .Q_t(n4406_t)
  );


  nnd2s3
  U3309
  (
    .DIN1(n3178),
    .DIN1_t(n3178_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4404),
    .Q_t(n4404_t)
  );


  xor2s3
  U3310
  (
    .DIN1(n4409),
    .DIN1_t(n4409_t),
    .DIN2(n4410),
    .DIN2_t(n4410_t),
    .Q(n3178),
    .Q_t(n3178_t)
  );


  xor2s3
  U3311
  (
    .DIN1(n6013),
    .DIN1_t(n6013_t),
    .DIN2(n4411),
    .DIN2_t(n4411_t),
    .Q(n4410),
    .Q_t(n4410_t)
  );


  xor2s3
  U3312
  (
    .DIN1(n6011),
    .DIN1_t(n6011_t),
    .DIN2(n6012),
    .DIN2_t(n6012_t),
    .Q(n4411),
    .Q_t(n4411_t)
  );


  xor2s3
  U3313
  (
    .DIN1(n6014),
    .DIN1_t(n6014_t),
    .DIN2(n6693),
    .DIN2_t(n6693_t),
    .Q(n4409),
    .Q_t(n4409_t)
  );


  nnd2s3
  U3314
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2229),
    .DIN2_t(n2229_t),
    .Q(n4403),
    .Q_t(n4403_t)
  );


  nnd2s3
  U3315
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2188),
    .DIN2_t(n2188_t),
    .Q(n4402),
    .Q_t(n4402_t)
  );


  nnd4s2
  U3316
  (
    .DIN1(n4412),
    .DIN1_t(n4412_t),
    .DIN2(n4413),
    .DIN2_t(n4413_t),
    .DIN3(n4414),
    .DIN3_t(n4414_t),
    .DIN4(n4415),
    .DIN4_t(n4415_t),
    .Q(WX1957),
    .Q_t(WX1957_t)
  );


  nnd2s3
  U3317
  (
    .DIN1(n4118),
    .DIN1_t(n4118_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4415),
    .Q_t(n4415_t)
  );


  xor2s3
  U3318
  (
    .DIN1(n4416),
    .DIN1_t(n4416_t),
    .DIN2(n4417),
    .DIN2_t(n4417_t),
    .Q(n4118),
    .Q_t(n4118_t)
  );


  xor2s3
  U3319
  (
    .DIN1(n6018),
    .DIN1_t(n6018_t),
    .DIN2(n4418),
    .DIN2_t(n4418_t),
    .Q(n4417),
    .Q_t(n4417_t)
  );


  xor2s3
  U3320
  (
    .DIN1(n6016),
    .DIN1_t(n6016_t),
    .DIN2(n6017),
    .DIN2_t(n6017_t),
    .Q(n4418),
    .Q_t(n4418_t)
  );


  xor2s3
  U3321
  (
    .DIN1(n6019),
    .DIN1_t(n6019_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4416),
    .Q_t(n4416_t)
  );


  nnd2s3
  U3322
  (
    .DIN1(n3184),
    .DIN1_t(n3184_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4414),
    .Q_t(n4414_t)
  );


  xor2s3
  U3323
  (
    .DIN1(n4419),
    .DIN1_t(n4419_t),
    .DIN2(n4420),
    .DIN2_t(n4420_t),
    .Q(n3184),
    .Q_t(n3184_t)
  );


  xor2s3
  U3324
  (
    .DIN1(n6022),
    .DIN1_t(n6022_t),
    .DIN2(n4421),
    .DIN2_t(n4421_t),
    .Q(n4420),
    .Q_t(n4420_t)
  );


  xor2s3
  U3325
  (
    .DIN1(n6020),
    .DIN1_t(n6020_t),
    .DIN2(n6021),
    .DIN2_t(n6021_t),
    .Q(n4421),
    .Q_t(n4421_t)
  );


  xor2s3
  U3326
  (
    .DIN1(n6023),
    .DIN1_t(n6023_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4419),
    .Q_t(n4419_t)
  );


  nnd2s3
  U3327
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2230),
    .DIN2_t(n2230_t),
    .Q(n4413),
    .Q_t(n4413_t)
  );


  nnd2s3
  U3328
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2187),
    .DIN2_t(n2187_t),
    .Q(n4412),
    .Q_t(n4412_t)
  );


  nnd4s2
  U3329
  (
    .DIN1(n4422),
    .DIN1_t(n4422_t),
    .DIN2(n4423),
    .DIN2_t(n4423_t),
    .DIN3(n4424),
    .DIN3_t(n4424_t),
    .DIN4(n4425),
    .DIN4_t(n4425_t),
    .Q(WX1955),
    .Q_t(WX1955_t)
  );


  nnd2s3
  U3330
  (
    .DIN1(n4126),
    .DIN1_t(n4126_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4425),
    .Q_t(n4425_t)
  );


  xor2s3
  U3331
  (
    .DIN1(n4426),
    .DIN1_t(n4426_t),
    .DIN2(n4427),
    .DIN2_t(n4427_t),
    .Q(n4126),
    .Q_t(n4126_t)
  );


  xor2s3
  U3332
  (
    .DIN1(n6027),
    .DIN1_t(n6027_t),
    .DIN2(n4428),
    .DIN2_t(n4428_t),
    .Q(n4427),
    .Q_t(n4427_t)
  );


  xor2s3
  U3333
  (
    .DIN1(n6025),
    .DIN1_t(n6025_t),
    .DIN2(n6026),
    .DIN2_t(n6026_t),
    .Q(n4428),
    .Q_t(n4428_t)
  );


  xor2s3
  U3334
  (
    .DIN1(n6028),
    .DIN1_t(n6028_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4426),
    .Q_t(n4426_t)
  );


  nnd2s3
  U3335
  (
    .DIN1(n3190),
    .DIN1_t(n3190_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4424),
    .Q_t(n4424_t)
  );


  xor2s3
  U3336
  (
    .DIN1(n4429),
    .DIN1_t(n4429_t),
    .DIN2(n4430),
    .DIN2_t(n4430_t),
    .Q(n3190),
    .Q_t(n3190_t)
  );


  xor2s3
  U3337
  (
    .DIN1(n6031),
    .DIN1_t(n6031_t),
    .DIN2(n4431),
    .DIN2_t(n4431_t),
    .Q(n4430),
    .Q_t(n4430_t)
  );


  xor2s3
  U3338
  (
    .DIN1(n6029),
    .DIN1_t(n6029_t),
    .DIN2(n6030),
    .DIN2_t(n6030_t),
    .Q(n4431),
    .Q_t(n4431_t)
  );


  xor2s3
  U3339
  (
    .DIN1(n6032),
    .DIN1_t(n6032_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4429),
    .Q_t(n4429_t)
  );


  nnd2s3
  U3340
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2231),
    .DIN2_t(n2231_t),
    .Q(n4423),
    .Q_t(n4423_t)
  );


  nnd2s3
  U3341
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2186),
    .DIN2_t(n2186_t),
    .Q(n4422),
    .Q_t(n4422_t)
  );


  nnd4s2
  U3342
  (
    .DIN1(n4432),
    .DIN1_t(n4432_t),
    .DIN2(n4433),
    .DIN2_t(n4433_t),
    .DIN3(n4434),
    .DIN3_t(n4434_t),
    .DIN4(n4435),
    .DIN4_t(n4435_t),
    .Q(WX1953),
    .Q_t(WX1953_t)
  );


  nnd2s3
  U3343
  (
    .DIN1(n4134),
    .DIN1_t(n4134_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4435),
    .Q_t(n4435_t)
  );


  xor2s3
  U3344
  (
    .DIN1(n4436),
    .DIN1_t(n4436_t),
    .DIN2(n4437),
    .DIN2_t(n4437_t),
    .Q(n4134),
    .Q_t(n4134_t)
  );


  xor2s3
  U3345
  (
    .DIN1(n6036),
    .DIN1_t(n6036_t),
    .DIN2(n4438),
    .DIN2_t(n4438_t),
    .Q(n4437),
    .Q_t(n4437_t)
  );


  xor2s3
  U3346
  (
    .DIN1(n6034),
    .DIN1_t(n6034_t),
    .DIN2(n6035),
    .DIN2_t(n6035_t),
    .Q(n4438),
    .Q_t(n4438_t)
  );


  xor2s3
  U3347
  (
    .DIN1(n6037),
    .DIN1_t(n6037_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4436),
    .Q_t(n4436_t)
  );


  nnd2s3
  U3348
  (
    .DIN1(n3196),
    .DIN1_t(n3196_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4434),
    .Q_t(n4434_t)
  );


  xor2s3
  U3349
  (
    .DIN1(n4439),
    .DIN1_t(n4439_t),
    .DIN2(n4440),
    .DIN2_t(n4440_t),
    .Q(n3196),
    .Q_t(n3196_t)
  );


  xor2s3
  U3350
  (
    .DIN1(n6040),
    .DIN1_t(n6040_t),
    .DIN2(n4441),
    .DIN2_t(n4441_t),
    .Q(n4440),
    .Q_t(n4440_t)
  );


  xor2s3
  U3351
  (
    .DIN1(n6038),
    .DIN1_t(n6038_t),
    .DIN2(n6039),
    .DIN2_t(n6039_t),
    .Q(n4441),
    .Q_t(n4441_t)
  );


  xor2s3
  U3352
  (
    .DIN1(n6041),
    .DIN1_t(n6041_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4439),
    .Q_t(n4439_t)
  );


  nnd2s3
  U3353
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2232),
    .DIN2_t(n2232_t),
    .Q(n4433),
    .Q_t(n4433_t)
  );


  nnd2s3
  U3354
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2185),
    .DIN2_t(n2185_t),
    .Q(n4432),
    .Q_t(n4432_t)
  );


  nnd4s2
  U3355
  (
    .DIN1(n4442),
    .DIN1_t(n4442_t),
    .DIN2(n4443),
    .DIN2_t(n4443_t),
    .DIN3(n4444),
    .DIN3_t(n4444_t),
    .DIN4(n4445),
    .DIN4_t(n4445_t),
    .Q(WX1951),
    .Q_t(WX1951_t)
  );


  nnd2s3
  U3356
  (
    .DIN1(n4142),
    .DIN1_t(n4142_t),
    .DIN2(n6639),
    .DIN2_t(n6639_t),
    .Q(n4445),
    .Q_t(n4445_t)
  );


  xor2s3
  U3357
  (
    .DIN1(n4446),
    .DIN1_t(n4446_t),
    .DIN2(n4447),
    .DIN2_t(n4447_t),
    .Q(n4142),
    .Q_t(n4142_t)
  );


  xor2s3
  U3358
  (
    .DIN1(n6045),
    .DIN1_t(n6045_t),
    .DIN2(n4448),
    .DIN2_t(n4448_t),
    .Q(n4447),
    .Q_t(n4447_t)
  );


  xor2s3
  U3359
  (
    .DIN1(n6043),
    .DIN1_t(n6043_t),
    .DIN2(n6044),
    .DIN2_t(n6044_t),
    .Q(n4448),
    .Q_t(n4448_t)
  );


  xor2s3
  U3360
  (
    .DIN1(n6046),
    .DIN1_t(n6046_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4446),
    .Q_t(n4446_t)
  );


  nnd2s3
  U3361
  (
    .DIN1(n3202),
    .DIN1_t(n3202_t),
    .DIN2(n6670),
    .DIN2_t(n6670_t),
    .Q(n4444),
    .Q_t(n4444_t)
  );


  xor2s3
  U3362
  (
    .DIN1(n4449),
    .DIN1_t(n4449_t),
    .DIN2(n4450),
    .DIN2_t(n4450_t),
    .Q(n3202),
    .Q_t(n3202_t)
  );


  xor2s3
  U3363
  (
    .DIN1(n6049),
    .DIN1_t(n6049_t),
    .DIN2(n4451),
    .DIN2_t(n4451_t),
    .Q(n4450),
    .Q_t(n4450_t)
  );


  xor2s3
  U3364
  (
    .DIN1(n6047),
    .DIN1_t(n6047_t),
    .DIN2(n6048),
    .DIN2_t(n6048_t),
    .Q(n4451),
    .Q_t(n4451_t)
  );


  xor2s3
  U3365
  (
    .DIN1(n6050),
    .DIN1_t(n6050_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4449),
    .Q_t(n4449_t)
  );


  nnd2s3
  U3366
  (
    .DIN1(n6597),
    .DIN1_t(n6597_t),
    .DIN2(n2233),
    .DIN2_t(n2233_t),
    .Q(n4443),
    .Q_t(n4443_t)
  );


  nnd2s3
  U3367
  (
    .DIN1(n6566),
    .DIN1_t(n6566_t),
    .DIN2(n2184),
    .DIN2_t(n2184_t),
    .Q(n4442),
    .Q_t(n4442_t)
  );


  nnd4s2
  U3368
  (
    .DIN1(n4452),
    .DIN1_t(n4452_t),
    .DIN2(n4453),
    .DIN2_t(n4453_t),
    .DIN3(n4454),
    .DIN3_t(n4454_t),
    .DIN4(n4455),
    .DIN4_t(n4455_t),
    .Q(WX1949),
    .Q_t(WX1949_t)
  );


  nnd2s3
  U3369
  (
    .DIN1(n4150),
    .DIN1_t(n4150_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4455),
    .Q_t(n4455_t)
  );


  xor2s3
  U3370
  (
    .DIN1(n4456),
    .DIN1_t(n4456_t),
    .DIN2(n4457),
    .DIN2_t(n4457_t),
    .Q(n4150),
    .Q_t(n4150_t)
  );


  xor2s3
  U3371
  (
    .DIN1(n6054),
    .DIN1_t(n6054_t),
    .DIN2(n4458),
    .DIN2_t(n4458_t),
    .Q(n4457),
    .Q_t(n4457_t)
  );


  xor2s3
  U3372
  (
    .DIN1(n6052),
    .DIN1_t(n6052_t),
    .DIN2(n6053),
    .DIN2_t(n6053_t),
    .Q(n4458),
    .Q_t(n4458_t)
  );


  xor2s3
  U3373
  (
    .DIN1(n6055),
    .DIN1_t(n6055_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4456),
    .Q_t(n4456_t)
  );


  nnd2s3
  U3374
  (
    .DIN1(n3336),
    .DIN1_t(n3336_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4454),
    .Q_t(n4454_t)
  );


  xor2s3
  U3375
  (
    .DIN1(n4459),
    .DIN1_t(n4459_t),
    .DIN2(n4460),
    .DIN2_t(n4460_t),
    .Q(n3336),
    .Q_t(n3336_t)
  );


  xor2s3
  U3376
  (
    .DIN1(n6058),
    .DIN1_t(n6058_t),
    .DIN2(n4461),
    .DIN2_t(n4461_t),
    .Q(n4460),
    .Q_t(n4460_t)
  );


  xor2s3
  U3377
  (
    .DIN1(n6056),
    .DIN1_t(n6056_t),
    .DIN2(n6057),
    .DIN2_t(n6057_t),
    .Q(n4461),
    .Q_t(n4461_t)
  );


  xor2s3
  U3378
  (
    .DIN1(n6059),
    .DIN1_t(n6059_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4459),
    .Q_t(n4459_t)
  );


  nnd2s3
  U3379
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n2234),
    .DIN2_t(n2234_t),
    .Q(n4453),
    .Q_t(n4453_t)
  );


  nnd2s3
  U3380
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n2183),
    .DIN2_t(n2183_t),
    .Q(n4452),
    .Q_t(n4452_t)
  );


  nnd4s2
  U3381
  (
    .DIN1(n4462),
    .DIN1_t(n4462_t),
    .DIN2(n4463),
    .DIN2_t(n4463_t),
    .DIN3(n4464),
    .DIN3_t(n4464_t),
    .DIN4(n4465),
    .DIN4_t(n4465_t),
    .Q(WX1947),
    .Q_t(WX1947_t)
  );


  nnd2s3
  U3382
  (
    .DIN1(n4158),
    .DIN1_t(n4158_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4465),
    .Q_t(n4465_t)
  );


  xor2s3
  U3383
  (
    .DIN1(n4466),
    .DIN1_t(n4466_t),
    .DIN2(n4467),
    .DIN2_t(n4467_t),
    .Q(n4158),
    .Q_t(n4158_t)
  );


  xor2s3
  U3384
  (
    .DIN1(n6063),
    .DIN1_t(n6063_t),
    .DIN2(n4468),
    .DIN2_t(n4468_t),
    .Q(n4467),
    .Q_t(n4467_t)
  );


  xor2s3
  U3385
  (
    .DIN1(n6061),
    .DIN1_t(n6061_t),
    .DIN2(n6062),
    .DIN2_t(n6062_t),
    .Q(n4468),
    .Q_t(n4468_t)
  );


  xor2s3
  U3386
  (
    .DIN1(n6064),
    .DIN1_t(n6064_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4466),
    .Q_t(n4466_t)
  );


  nnd2s3
  U3387
  (
    .DIN1(n3342),
    .DIN1_t(n3342_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4464),
    .Q_t(n4464_t)
  );


  xor2s3
  U3388
  (
    .DIN1(n4469),
    .DIN1_t(n4469_t),
    .DIN2(n4470),
    .DIN2_t(n4470_t),
    .Q(n3342),
    .Q_t(n3342_t)
  );


  xor2s3
  U3389
  (
    .DIN1(n6067),
    .DIN1_t(n6067_t),
    .DIN2(n4471),
    .DIN2_t(n4471_t),
    .Q(n4470),
    .Q_t(n4470_t)
  );


  xor2s3
  U3390
  (
    .DIN1(n6065),
    .DIN1_t(n6065_t),
    .DIN2(n6066),
    .DIN2_t(n6066_t),
    .Q(n4471),
    .Q_t(n4471_t)
  );


  xor2s3
  U3391
  (
    .DIN1(n6068),
    .DIN1_t(n6068_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4469),
    .Q_t(n4469_t)
  );


  nnd2s3
  U3392
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n2235),
    .DIN2_t(n2235_t),
    .Q(n4463),
    .Q_t(n4463_t)
  );


  nnd2s3
  U3393
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n2182),
    .DIN2_t(n2182_t),
    .Q(n4462),
    .Q_t(n4462_t)
  );


  nnd4s2
  U3394
  (
    .DIN1(n4472),
    .DIN1_t(n4472_t),
    .DIN2(n4473),
    .DIN2_t(n4473_t),
    .DIN3(n4474),
    .DIN3_t(n4474_t),
    .DIN4(n4475),
    .DIN4_t(n4475_t),
    .Q(WX1945),
    .Q_t(WX1945_t)
  );


  nnd2s3
  U3395
  (
    .DIN1(n4166),
    .DIN1_t(n4166_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4475),
    .Q_t(n4475_t)
  );


  xor2s3
  U3396
  (
    .DIN1(n4476),
    .DIN1_t(n4476_t),
    .DIN2(n4477),
    .DIN2_t(n4477_t),
    .Q(n4166),
    .Q_t(n4166_t)
  );


  xor2s3
  U3397
  (
    .DIN1(n6072),
    .DIN1_t(n6072_t),
    .DIN2(n4478),
    .DIN2_t(n4478_t),
    .Q(n4477),
    .Q_t(n4477_t)
  );


  xor2s3
  U3398
  (
    .DIN1(n6070),
    .DIN1_t(n6070_t),
    .DIN2(n6071),
    .DIN2_t(n6071_t),
    .Q(n4478),
    .Q_t(n4478_t)
  );


  xor2s3
  U3399
  (
    .DIN1(n6073),
    .DIN1_t(n6073_t),
    .DIN2(n6694),
    .DIN2_t(n6694_t),
    .Q(n4476),
    .Q_t(n4476_t)
  );


  nnd2s3
  U3400
  (
    .DIN1(n3348),
    .DIN1_t(n3348_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4474),
    .Q_t(n4474_t)
  );


  xor2s3
  U3401
  (
    .DIN1(n4479),
    .DIN1_t(n4479_t),
    .DIN2(n4480),
    .DIN2_t(n4480_t),
    .Q(n3348),
    .Q_t(n3348_t)
  );


  xor2s3
  U3402
  (
    .DIN1(n6076),
    .DIN1_t(n6076_t),
    .DIN2(n4481),
    .DIN2_t(n4481_t),
    .Q(n4480),
    .Q_t(n4480_t)
  );


  xor2s3
  U3403
  (
    .DIN1(n6074),
    .DIN1_t(n6074_t),
    .DIN2(n6075),
    .DIN2_t(n6075_t),
    .Q(n4481),
    .Q_t(n4481_t)
  );


  xor2s3
  U3404
  (
    .DIN1(n6077),
    .DIN1_t(n6077_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4479),
    .Q_t(n4479_t)
  );


  nnd2s3
  U3405
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n2236),
    .DIN2_t(n2236_t),
    .Q(n4473),
    .Q_t(n4473_t)
  );


  nnd2s3
  U3406
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n2181),
    .DIN2_t(n2181_t),
    .Q(n4472),
    .Q_t(n4472_t)
  );


  nnd4s2
  U3407
  (
    .DIN1(n4482),
    .DIN1_t(n4482_t),
    .DIN2(n4483),
    .DIN2_t(n4483_t),
    .DIN3(n4484),
    .DIN3_t(n4484_t),
    .DIN4(n4485),
    .DIN4_t(n4485_t),
    .Q(WX1943),
    .Q_t(WX1943_t)
  );


  nnd2s3
  U3408
  (
    .DIN1(n4174),
    .DIN1_t(n4174_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4485),
    .Q_t(n4485_t)
  );


  xor2s3
  U3409
  (
    .DIN1(n4486),
    .DIN1_t(n4486_t),
    .DIN2(n4487),
    .DIN2_t(n4487_t),
    .Q(n4174),
    .Q_t(n4174_t)
  );


  xor2s3
  U3410
  (
    .DIN1(n6081),
    .DIN1_t(n6081_t),
    .DIN2(n4488),
    .DIN2_t(n4488_t),
    .Q(n4487),
    .Q_t(n4487_t)
  );


  xor2s3
  U3411
  (
    .DIN1(n6079),
    .DIN1_t(n6079_t),
    .DIN2(n6080),
    .DIN2_t(n6080_t),
    .Q(n4488),
    .Q_t(n4488_t)
  );


  xor2s3
  U3412
  (
    .DIN1(n6082),
    .DIN1_t(n6082_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4486),
    .Q_t(n4486_t)
  );


  nnd2s3
  U3413
  (
    .DIN1(n3354),
    .DIN1_t(n3354_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4484),
    .Q_t(n4484_t)
  );


  xor2s3
  U3414
  (
    .DIN1(n4489),
    .DIN1_t(n4489_t),
    .DIN2(n4490),
    .DIN2_t(n4490_t),
    .Q(n3354),
    .Q_t(n3354_t)
  );


  xor2s3
  U3415
  (
    .DIN1(n6085),
    .DIN1_t(n6085_t),
    .DIN2(n4491),
    .DIN2_t(n4491_t),
    .Q(n4490),
    .Q_t(n4490_t)
  );


  xor2s3
  U3416
  (
    .DIN1(n6083),
    .DIN1_t(n6083_t),
    .DIN2(n6084),
    .DIN2_t(n6084_t),
    .Q(n4491),
    .Q_t(n4491_t)
  );


  xor2s3
  U3417
  (
    .DIN1(n6086),
    .DIN1_t(n6086_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4489),
    .Q_t(n4489_t)
  );


  nnd2s3
  U3418
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n2237),
    .DIN2_t(n2237_t),
    .Q(n4483),
    .Q_t(n4483_t)
  );


  nnd2s3
  U3419
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n2180),
    .DIN2_t(n2180_t),
    .Q(n4482),
    .Q_t(n4482_t)
  );


  nnd4s2
  U3420
  (
    .DIN1(n4492),
    .DIN1_t(n4492_t),
    .DIN2(n4493),
    .DIN2_t(n4493_t),
    .DIN3(n4494),
    .DIN3_t(n4494_t),
    .DIN4(n4495),
    .DIN4_t(n4495_t),
    .Q(WX1941),
    .Q_t(WX1941_t)
  );


  nnd2s3
  U3421
  (
    .DIN1(n4182),
    .DIN1_t(n4182_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4495),
    .Q_t(n4495_t)
  );


  xor2s3
  U3422
  (
    .DIN1(n4496),
    .DIN1_t(n4496_t),
    .DIN2(n4497),
    .DIN2_t(n4497_t),
    .Q(n4182),
    .Q_t(n4182_t)
  );


  xor2s3
  U3423
  (
    .DIN1(n6090),
    .DIN1_t(n6090_t),
    .DIN2(n4498),
    .DIN2_t(n4498_t),
    .Q(n4497),
    .Q_t(n4497_t)
  );


  xor2s3
  U3424
  (
    .DIN1(n6088),
    .DIN1_t(n6088_t),
    .DIN2(n6089),
    .DIN2_t(n6089_t),
    .Q(n4498),
    .Q_t(n4498_t)
  );


  xor2s3
  U3425
  (
    .DIN1(n6091),
    .DIN1_t(n6091_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4496),
    .Q_t(n4496_t)
  );


  nnd2s3
  U3426
  (
    .DIN1(n3370),
    .DIN1_t(n3370_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4494),
    .Q_t(n4494_t)
  );


  xor2s3
  U3427
  (
    .DIN1(n4499),
    .DIN1_t(n4499_t),
    .DIN2(n4500),
    .DIN2_t(n4500_t),
    .Q(n3370),
    .Q_t(n3370_t)
  );


  xor2s3
  U3428
  (
    .DIN1(n6094),
    .DIN1_t(n6094_t),
    .DIN2(n4501),
    .DIN2_t(n4501_t),
    .Q(n4500),
    .Q_t(n4500_t)
  );


  xor2s3
  U3429
  (
    .DIN1(n6092),
    .DIN1_t(n6092_t),
    .DIN2(n6093),
    .DIN2_t(n6093_t),
    .Q(n4501),
    .Q_t(n4501_t)
  );


  xor2s3
  U3430
  (
    .DIN1(n6095),
    .DIN1_t(n6095_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4499),
    .Q_t(n4499_t)
  );


  nnd2s3
  U3431
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n2238),
    .DIN2_t(n2238_t),
    .Q(n4493),
    .Q_t(n4493_t)
  );


  nnd2s3
  U3432
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n2179),
    .DIN2_t(n2179_t),
    .Q(n4492),
    .Q_t(n4492_t)
  );


  nnd4s2
  U3433
  (
    .DIN1(n4502),
    .DIN1_t(n4502_t),
    .DIN2(n4503),
    .DIN2_t(n4503_t),
    .DIN3(n4504),
    .DIN3_t(n4504_t),
    .DIN4(n4505),
    .DIN4_t(n4505_t),
    .Q(WX1939),
    .Q_t(WX1939_t)
  );


  nnd2s3
  U3434
  (
    .DIN1(n4190),
    .DIN1_t(n4190_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4505),
    .Q_t(n4505_t)
  );


  xor2s3
  U3435
  (
    .DIN1(n4506),
    .DIN1_t(n4506_t),
    .DIN2(n4507),
    .DIN2_t(n4507_t),
    .Q(n4190),
    .Q_t(n4190_t)
  );


  xor2s3
  U3436
  (
    .DIN1(n6099),
    .DIN1_t(n6099_t),
    .DIN2(n4508),
    .DIN2_t(n4508_t),
    .Q(n4507),
    .Q_t(n4507_t)
  );


  xor2s3
  U3437
  (
    .DIN1(n6097),
    .DIN1_t(n6097_t),
    .DIN2(n6098),
    .DIN2_t(n6098_t),
    .Q(n4508),
    .Q_t(n4508_t)
  );


  xor2s3
  U3438
  (
    .DIN1(n6100),
    .DIN1_t(n6100_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4506),
    .Q_t(n4506_t)
  );


  nnd2s3
  U3439
  (
    .DIN1(n3387),
    .DIN1_t(n3387_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4504),
    .Q_t(n4504_t)
  );


  xor2s3
  U3440
  (
    .DIN1(n4509),
    .DIN1_t(n4509_t),
    .DIN2(n4510),
    .DIN2_t(n4510_t),
    .Q(n3387),
    .Q_t(n3387_t)
  );


  xor2s3
  U3441
  (
    .DIN1(n6103),
    .DIN1_t(n6103_t),
    .DIN2(n4511),
    .DIN2_t(n4511_t),
    .Q(n4510),
    .Q_t(n4510_t)
  );


  xor2s3
  U3442
  (
    .DIN1(n6101),
    .DIN1_t(n6101_t),
    .DIN2(n6102),
    .DIN2_t(n6102_t),
    .Q(n4511),
    .Q_t(n4511_t)
  );


  xor2s3
  U3443
  (
    .DIN1(n6104),
    .DIN1_t(n6104_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4509),
    .Q_t(n4509_t)
  );


  nnd2s3
  U3444
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n2239),
    .DIN2_t(n2239_t),
    .Q(n4503),
    .Q_t(n4503_t)
  );


  nnd2s3
  U3445
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n2178),
    .DIN2_t(n2178_t),
    .Q(n4502),
    .Q_t(n4502_t)
  );


  nnd4s2
  U3446
  (
    .DIN1(n4512),
    .DIN1_t(n4512_t),
    .DIN2(n4513),
    .DIN2_t(n4513_t),
    .DIN3(n4514),
    .DIN3_t(n4514_t),
    .DIN4(n4515),
    .DIN4_t(n4515_t),
    .Q(WX1937),
    .Q_t(WX1937_t)
  );


  nnd2s3
  U3447
  (
    .DIN1(n4198),
    .DIN1_t(n4198_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4515),
    .Q_t(n4515_t)
  );


  xor2s3
  U3448
  (
    .DIN1(n4516),
    .DIN1_t(n4516_t),
    .DIN2(n4517),
    .DIN2_t(n4517_t),
    .Q(n4198),
    .Q_t(n4198_t)
  );


  xor2s3
  U3449
  (
    .DIN1(n6108),
    .DIN1_t(n6108_t),
    .DIN2(n4518),
    .DIN2_t(n4518_t),
    .Q(n4517),
    .Q_t(n4517_t)
  );


  xor2s3
  U3450
  (
    .DIN1(n6106),
    .DIN1_t(n6106_t),
    .DIN2(n6107),
    .DIN2_t(n6107_t),
    .Q(n4518),
    .Q_t(n4518_t)
  );


  xor2s3
  U3451
  (
    .DIN1(n6109),
    .DIN1_t(n6109_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4516),
    .Q_t(n4516_t)
  );


  nnd2s3
  U3452
  (
    .DIN1(n3405),
    .DIN1_t(n3405_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4514),
    .Q_t(n4514_t)
  );


  xor2s3
  U3453
  (
    .DIN1(n4519),
    .DIN1_t(n4519_t),
    .DIN2(n4520),
    .DIN2_t(n4520_t),
    .Q(n3405),
    .Q_t(n3405_t)
  );


  xor2s3
  U3454
  (
    .DIN1(n6112),
    .DIN1_t(n6112_t),
    .DIN2(n4521),
    .DIN2_t(n4521_t),
    .Q(n4520),
    .Q_t(n4520_t)
  );


  xor2s3
  U3455
  (
    .DIN1(n6110),
    .DIN1_t(n6110_t),
    .DIN2(n6111),
    .DIN2_t(n6111_t),
    .Q(n4521),
    .Q_t(n4521_t)
  );


  xor2s3
  U3456
  (
    .DIN1(n6113),
    .DIN1_t(n6113_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4519),
    .Q_t(n4519_t)
  );


  nnd2s3
  U3457
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n2240),
    .DIN2_t(n2240_t),
    .Q(n4513),
    .Q_t(n4513_t)
  );


  nnd2s3
  U3458
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n2177),
    .DIN2_t(n2177_t),
    .Q(n4512),
    .Q_t(n4512_t)
  );


  nor2s3
  U3459
  (
    .DIN1(n6803),
    .DIN1_t(n6803_t),
    .DIN2(n2240),
    .DIN2_t(n2240_t),
    .Q(WX1839),
    .Q_t(WX1839_t)
  );


  nor2s3
  U3460
  (
    .DIN1(n6116),
    .DIN1_t(n6116_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX1837),
    .Q_t(WX1837_t)
  );


  nor2s3
  U3461
  (
    .DIN1(n6117),
    .DIN1_t(n6117_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX1835),
    .Q_t(WX1835_t)
  );


  nor2s3
  U3462
  (
    .DIN1(n6118),
    .DIN1_t(n6118_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX1833),
    .Q_t(WX1833_t)
  );


  nor2s3
  U3463
  (
    .DIN1(n6119),
    .DIN1_t(n6119_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX1831),
    .Q_t(WX1831_t)
  );


  nor2s3
  U3464
  (
    .DIN1(n6120),
    .DIN1_t(n6120_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX1829),
    .Q_t(WX1829_t)
  );


  nor2s3
  U3465
  (
    .DIN1(n6121),
    .DIN1_t(n6121_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX1827),
    .Q_t(WX1827_t)
  );


  nor2s3
  U3466
  (
    .DIN1(n6122),
    .DIN1_t(n6122_t),
    .DIN2(n6757),
    .DIN2_t(n6757_t),
    .Q(WX1825),
    .Q_t(WX1825_t)
  );


  nor2s3
  U3467
  (
    .DIN1(n6123),
    .DIN1_t(n6123_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX1823),
    .Q_t(WX1823_t)
  );


  nor2s3
  U3468
  (
    .DIN1(n6124),
    .DIN1_t(n6124_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX1821),
    .Q_t(WX1821_t)
  );


  nor2s3
  U3469
  (
    .DIN1(n6125),
    .DIN1_t(n6125_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX1819),
    .Q_t(WX1819_t)
  );


  nor2s3
  U3470
  (
    .DIN1(n6126),
    .DIN1_t(n6126_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX1817),
    .Q_t(WX1817_t)
  );


  nor2s3
  U3471
  (
    .DIN1(n6127),
    .DIN1_t(n6127_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX1815),
    .Q_t(WX1815_t)
  );


  nor2s3
  U3472
  (
    .DIN1(n6128),
    .DIN1_t(n6128_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX1813),
    .Q_t(WX1813_t)
  );


  nor2s3
  U3473
  (
    .DIN1(n6129),
    .DIN1_t(n6129_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX1811),
    .Q_t(WX1811_t)
  );


  nor2s3
  U3474
  (
    .DIN1(n6130),
    .DIN1_t(n6130_t),
    .DIN2(n6756),
    .DIN2_t(n6756_t),
    .Q(WX1809),
    .Q_t(WX1809_t)
  );


  nor2s3
  U3475
  (
    .DIN1(n6131),
    .DIN1_t(n6131_t),
    .DIN2(n6761),
    .DIN2_t(n6761_t),
    .Q(WX1807),
    .Q_t(WX1807_t)
  );


  nor2s3
  U3476
  (
    .DIN1(n6132),
    .DIN1_t(n6132_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1805),
    .Q_t(WX1805_t)
  );


  nor2s3
  U3477
  (
    .DIN1(n6133),
    .DIN1_t(n6133_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1803),
    .Q_t(WX1803_t)
  );


  nor2s3
  U3478
  (
    .DIN1(n6134),
    .DIN1_t(n6134_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1801),
    .Q_t(WX1801_t)
  );


  nor2s3
  U3479
  (
    .DIN1(n6135),
    .DIN1_t(n6135_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1799),
    .Q_t(WX1799_t)
  );


  nor2s3
  U3480
  (
    .DIN1(n6136),
    .DIN1_t(n6136_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1797),
    .Q_t(WX1797_t)
  );


  nor2s3
  U3481
  (
    .DIN1(n6137),
    .DIN1_t(n6137_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1795),
    .Q_t(WX1795_t)
  );


  nor2s3
  U3482
  (
    .DIN1(n6138),
    .DIN1_t(n6138_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1793),
    .Q_t(WX1793_t)
  );


  nor2s3
  U3483
  (
    .DIN1(n6139),
    .DIN1_t(n6139_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1791),
    .Q_t(WX1791_t)
  );


  nor2s3
  U3484
  (
    .DIN1(n6140),
    .DIN1_t(n6140_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1789),
    .Q_t(WX1789_t)
  );


  nor2s3
  U3485
  (
    .DIN1(n6141),
    .DIN1_t(n6141_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1787),
    .Q_t(WX1787_t)
  );


  nor2s3
  U3486
  (
    .DIN1(n6142),
    .DIN1_t(n6142_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1785),
    .Q_t(WX1785_t)
  );


  nor2s3
  U3487
  (
    .DIN1(n6143),
    .DIN1_t(n6143_t),
    .DIN2(n6775),
    .DIN2_t(n6775_t),
    .Q(WX1783),
    .Q_t(WX1783_t)
  );


  nor2s3
  U3488
  (
    .DIN1(n6144),
    .DIN1_t(n6144_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX1781),
    .Q_t(WX1781_t)
  );


  nor2s3
  U3489
  (
    .DIN1(n6145),
    .DIN1_t(n6145_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX1779),
    .Q_t(WX1779_t)
  );


  nor2s3
  U3490
  (
    .DIN1(n6146),
    .DIN1_t(n6146_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX1777),
    .Q_t(WX1777_t)
  );


  nor2s3
  U3491
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n4522),
    .DIN2_t(n4522_t),
    .Q(WX1326),
    .Q_t(WX1326_t)
  );


  xor2s3
  U3492
  (
    .DIN1(n6147),
    .DIN1_t(n6147_t),
    .DIN2(n6534),
    .DIN2_t(n6534_t),
    .Q(n4522),
    .Q_t(n4522_t)
  );


  nor2s3
  U3493
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n4523),
    .DIN2_t(n4523_t),
    .Q(WX1324),
    .Q_t(WX1324_t)
  );


  xor2s3
  U3494
  (
    .DIN1(n6148),
    .DIN1_t(n6148_t),
    .DIN2(n6474),
    .DIN2_t(n6474_t),
    .Q(n4523),
    .Q_t(n4523_t)
  );


  nor2s3
  U3495
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n4524),
    .DIN2_t(n4524_t),
    .Q(WX1322),
    .Q_t(WX1322_t)
  );


  xor2s3
  U3496
  (
    .DIN1(n6149),
    .DIN1_t(n6149_t),
    .DIN2(n6482),
    .DIN2_t(n6482_t),
    .Q(n4524),
    .Q_t(n4524_t)
  );


  nor2s3
  U3497
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n4525),
    .DIN2_t(n4525_t),
    .Q(WX1320),
    .Q_t(WX1320_t)
  );


  xor2s3
  U3498
  (
    .DIN1(n6150),
    .DIN1_t(n6150_t),
    .DIN2(n6483),
    .DIN2_t(n6483_t),
    .Q(n4525),
    .Q_t(n4525_t)
  );


  nor2s3
  U3499
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n4526),
    .DIN2_t(n4526_t),
    .Q(WX1318),
    .Q_t(WX1318_t)
  );


  xor2s3
  U3500
  (
    .DIN1(n6151),
    .DIN1_t(n6151_t),
    .DIN2(n6486),
    .DIN2_t(n6486_t),
    .Q(n4526),
    .Q_t(n4526_t)
  );


  nor2s3
  U3501
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n4527),
    .DIN2_t(n4527_t),
    .Q(WX1316),
    .Q_t(WX1316_t)
  );


  xor2s3
  U3502
  (
    .DIN1(n6152),
    .DIN1_t(n6152_t),
    .DIN2(n6492),
    .DIN2_t(n6492_t),
    .Q(n4527),
    .Q_t(n4527_t)
  );


  nor2s3
  U3503
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n4528),
    .DIN2_t(n4528_t),
    .Q(WX1314),
    .Q_t(WX1314_t)
  );


  xor2s3
  U3504
  (
    .DIN1(n6153),
    .DIN1_t(n6153_t),
    .DIN2(n6500),
    .DIN2_t(n6500_t),
    .Q(n4528),
    .Q_t(n4528_t)
  );


  nor2s3
  U3505
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n4529),
    .DIN2_t(n4529_t),
    .Q(WX1312),
    .Q_t(WX1312_t)
  );


  xor2s3
  U3506
  (
    .DIN1(n6154),
    .DIN1_t(n6154_t),
    .DIN2(n6501),
    .DIN2_t(n6501_t),
    .Q(n4529),
    .Q_t(n4529_t)
  );


  nor2s3
  U3507
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n4530),
    .DIN2_t(n4530_t),
    .Q(WX1310),
    .Q_t(WX1310_t)
  );


  xor2s3
  U3508
  (
    .DIN1(n6155),
    .DIN1_t(n6155_t),
    .DIN2(n6511),
    .DIN2_t(n6511_t),
    .Q(n4530),
    .Q_t(n4530_t)
  );


  nor2s3
  U3509
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n4531),
    .DIN2_t(n4531_t),
    .Q(WX1308),
    .Q_t(WX1308_t)
  );


  xor2s3
  U3510
  (
    .DIN1(n6156),
    .DIN1_t(n6156_t),
    .DIN2(n6516),
    .DIN2_t(n6516_t),
    .Q(n4531),
    .Q_t(n4531_t)
  );


  nor2s3
  U3511
  (
    .DIN1(n6805),
    .DIN1_t(n6805_t),
    .DIN2(n4532),
    .DIN2_t(n4532_t),
    .Q(WX1306),
    .Q_t(WX1306_t)
  );


  xor2s3
  U3512
  (
    .DIN1(n6157),
    .DIN1_t(n6157_t),
    .DIN2(n6517),
    .DIN2_t(n6517_t),
    .Q(n4532),
    .Q_t(n4532_t)
  );


  nor2s3
  U3513
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4533),
    .DIN2_t(n4533_t),
    .Q(WX1304),
    .Q_t(WX1304_t)
  );


  xor2s3
  U3514
  (
    .DIN1(n6158),
    .DIN1_t(n6158_t),
    .DIN2(n6522),
    .DIN2_t(n6522_t),
    .Q(n4533),
    .Q_t(n4533_t)
  );


  nor2s3
  U3515
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4534),
    .DIN2_t(n4534_t),
    .Q(WX1302),
    .Q_t(WX1302_t)
  );


  xor2s3
  U3516
  (
    .DIN1(n6159),
    .DIN1_t(n6159_t),
    .DIN2(n6477),
    .DIN2_t(n6477_t),
    .Q(n4534),
    .Q_t(n4534_t)
  );


  nor2s3
  U3517
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4535),
    .DIN2_t(n4535_t),
    .Q(WX1300),
    .Q_t(WX1300_t)
  );


  xor2s3
  U3518
  (
    .DIN1(n6160),
    .DIN1_t(n6160_t),
    .DIN2(n6491),
    .DIN2_t(n6491_t),
    .Q(n4535),
    .Q_t(n4535_t)
  );


  nor2s3
  U3519
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4536),
    .DIN2_t(n4536_t),
    .Q(WX1298),
    .Q_t(WX1298_t)
  );


  xor2s3
  U3520
  (
    .DIN1(n6161),
    .DIN1_t(n6161_t),
    .DIN2(n6495),
    .DIN2_t(n6495_t),
    .Q(n4536),
    .Q_t(n4536_t)
  );


  nor2s3
  U3521
  (
    .DIN1(n4537),
    .DIN1_t(n4537_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX1296),
    .Q_t(WX1296_t)
  );


  xnr2s3
  U3522
  (
    .DIN1(n6510),
    .DIN1_t(n6510_t),
    .DIN2(n4538),
    .DIN2_t(n4538_t),
    .Q(n4537),
    .Q_t(n4537_t)
  );


  xor2s3
  U3523
  (
    .DIN1(n6162),
    .DIN1_t(n6162_t),
    .DIN2(n6178),
    .DIN2_t(n6178_t),
    .Q(n4538),
    .Q_t(n4538_t)
  );


  nor2s3
  U3524
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4539),
    .DIN2_t(n4539_t),
    .Q(WX1294),
    .Q_t(WX1294_t)
  );


  xor2s3
  U3525
  (
    .DIN1(n6163),
    .DIN1_t(n6163_t),
    .DIN2(n6438),
    .DIN2_t(n6438_t),
    .Q(n4539),
    .Q_t(n4539_t)
  );


  nor2s3
  U3526
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4540),
    .DIN2_t(n4540_t),
    .Q(WX1292),
    .Q_t(WX1292_t)
  );


  xor2s3
  U3527
  (
    .DIN1(n6164),
    .DIN1_t(n6164_t),
    .DIN2(n6525),
    .DIN2_t(n6525_t),
    .Q(n4540),
    .Q_t(n4540_t)
  );


  nor2s3
  U3528
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4541),
    .DIN2_t(n4541_t),
    .Q(WX1290),
    .Q_t(WX1290_t)
  );


  xor2s3
  U3529
  (
    .DIN1(n6165),
    .DIN1_t(n6165_t),
    .DIN2(n6447),
    .DIN2_t(n6447_t),
    .Q(n4541),
    .Q_t(n4541_t)
  );


  nor2s3
  U3530
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4542),
    .DIN2_t(n4542_t),
    .Q(WX1288),
    .Q_t(WX1288_t)
  );


  xor2s3
  U3531
  (
    .DIN1(n6166),
    .DIN1_t(n6166_t),
    .DIN2(n6456),
    .DIN2_t(n6456_t),
    .Q(n4542),
    .Q_t(n4542_t)
  );


  nor2s3
  U3532
  (
    .DIN1(n4543),
    .DIN1_t(n4543_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX1286),
    .Q_t(WX1286_t)
  );


  xnr2s3
  U3533
  (
    .DIN1(n6444),
    .DIN1_t(n6444_t),
    .DIN2(n4544),
    .DIN2_t(n4544_t),
    .Q(n4543),
    .Q_t(n4543_t)
  );


  xor2s3
  U3534
  (
    .DIN1(n6167),
    .DIN1_t(n6167_t),
    .DIN2(n6178),
    .DIN2_t(n6178_t),
    .Q(n4544),
    .Q_t(n4544_t)
  );


  nor2s3
  U3535
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4545),
    .DIN2_t(n4545_t),
    .Q(WX1284),
    .Q_t(WX1284_t)
  );


  xor2s3
  U3536
  (
    .DIN1(n6168),
    .DIN1_t(n6168_t),
    .DIN2(n6450),
    .DIN2_t(n6450_t),
    .Q(n4545),
    .Q_t(n4545_t)
  );


  nor2s3
  U3537
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4546),
    .DIN2_t(n4546_t),
    .Q(WX1282),
    .Q_t(WX1282_t)
  );


  xor2s3
  U3538
  (
    .DIN1(n6169),
    .DIN1_t(n6169_t),
    .DIN2(n6506),
    .DIN2_t(n6506_t),
    .Q(n4546),
    .Q_t(n4546_t)
  );


  nor2s3
  U3539
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4547),
    .DIN2_t(n4547_t),
    .Q(WX1280),
    .Q_t(WX1280_t)
  );


  xor2s3
  U3540
  (
    .DIN1(n6170),
    .DIN1_t(n6170_t),
    .DIN2(n6453),
    .DIN2_t(n6453_t),
    .Q(n4547),
    .Q_t(n4547_t)
  );


  nor2s3
  U3541
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4548),
    .DIN2_t(n4548_t),
    .Q(WX1278),
    .Q_t(WX1278_t)
  );


  xor2s3
  U3542
  (
    .DIN1(n6171),
    .DIN1_t(n6171_t),
    .DIN2(n6465),
    .DIN2_t(n6465_t),
    .Q(n4548),
    .Q_t(n4548_t)
  );


  nor2s3
  U3543
  (
    .DIN1(n6806),
    .DIN1_t(n6806_t),
    .DIN2(n4549),
    .DIN2_t(n4549_t),
    .Q(WX1276),
    .Q_t(WX1276_t)
  );


  xor2s3
  U3544
  (
    .DIN1(n6172),
    .DIN1_t(n6172_t),
    .DIN2(n6441),
    .DIN2_t(n6441_t),
    .Q(n4549),
    .Q_t(n4549_t)
  );


  nor2s3
  U3545
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4550),
    .DIN2_t(n4550_t),
    .Q(WX1274),
    .Q_t(WX1274_t)
  );


  xor2s3
  U3546
  (
    .DIN1(n6173),
    .DIN1_t(n6173_t),
    .DIN2(n6459),
    .DIN2_t(n6459_t),
    .Q(n4550),
    .Q_t(n4550_t)
  );


  nor2s3
  U3547
  (
    .DIN1(n4551),
    .DIN1_t(n4551_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX1272),
    .Q_t(WX1272_t)
  );


  xnr2s3
  U3548
  (
    .DIN1(n6471),
    .DIN1_t(n6471_t),
    .DIN2(n4552),
    .DIN2_t(n4552_t),
    .Q(n4551),
    .Q_t(n4551_t)
  );


  xor2s3
  U3549
  (
    .DIN1(n6174),
    .DIN1_t(n6174_t),
    .DIN2(n6178),
    .DIN2_t(n6178_t),
    .Q(n4552),
    .Q_t(n4552_t)
  );


  nor2s3
  U3550
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4553),
    .DIN2_t(n4553_t),
    .Q(WX1270),
    .Q_t(WX1270_t)
  );


  xor2s3
  U3551
  (
    .DIN1(n6175),
    .DIN1_t(n6175_t),
    .DIN2(n6468),
    .DIN2_t(n6468_t),
    .Q(n4553),
    .Q_t(n4553_t)
  );


  nor2s3
  U3552
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4554),
    .DIN2_t(n4554_t),
    .Q(WX1268),
    .Q_t(WX1268_t)
  );


  xor2s3
  U3553
  (
    .DIN1(n6176),
    .DIN1_t(n6176_t),
    .DIN2(n6437),
    .DIN2_t(n6437_t),
    .Q(n4554),
    .Q_t(n4554_t)
  );


  nor2s3
  U3554
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4555),
    .DIN2_t(n4555_t),
    .Q(WX1266),
    .Q_t(WX1266_t)
  );


  xor2s3
  U3555
  (
    .DIN1(n6177),
    .DIN1_t(n6177_t),
    .DIN2(n6530),
    .DIN2_t(n6530_t),
    .Q(n4555),
    .Q_t(n4555_t)
  );


  nor2s3
  U3556
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4556),
    .DIN2_t(n4556_t),
    .Q(WX1264),
    .Q_t(WX1264_t)
  );


  xor2s3
  U3557
  (
    .DIN1(n6178),
    .DIN1_t(n6178_t),
    .DIN2(n6462),
    .DIN2_t(n6462_t),
    .Q(n4556),
    .Q_t(n4556_t)
  );


  nor2s3
  U3558
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4557),
    .DIN2_t(n4557_t),
    .Q(WX11670),
    .Q_t(WX11670_t)
  );


  xor2s3
  U3559
  (
    .DIN1(n6336),
    .DIN1_t(n6336_t),
    .DIN2(n6341),
    .DIN2_t(n6341_t),
    .Q(n4557),
    .Q_t(n4557_t)
  );


  nor2s3
  U3560
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4558),
    .DIN2_t(n4558_t),
    .Q(WX11668),
    .Q_t(WX11668_t)
  );


  xor2s3
  U3561
  (
    .DIN1(n6331),
    .DIN1_t(n6331_t),
    .DIN2(n6335),
    .DIN2_t(n6335_t),
    .Q(n4558),
    .Q_t(n4558_t)
  );


  nor2s3
  U3562
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4559),
    .DIN2_t(n4559_t),
    .Q(WX11666),
    .Q_t(WX11666_t)
  );


  xor2s3
  U3563
  (
    .DIN1(n6326),
    .DIN1_t(n6326_t),
    .DIN2(n6330),
    .DIN2_t(n6330_t),
    .Q(n4559),
    .Q_t(n4559_t)
  );


  nor2s3
  U3564
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4560),
    .DIN2_t(n4560_t),
    .Q(WX11664),
    .Q_t(WX11664_t)
  );


  xor2s3
  U3565
  (
    .DIN1(n6321),
    .DIN1_t(n6321_t),
    .DIN2(n6325),
    .DIN2_t(n6325_t),
    .Q(n4560),
    .Q_t(n4560_t)
  );


  nor2s3
  U3566
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4561),
    .DIN2_t(n4561_t),
    .Q(WX11662),
    .Q_t(WX11662_t)
  );


  xor2s3
  U3567
  (
    .DIN1(n6316),
    .DIN1_t(n6316_t),
    .DIN2(n6320),
    .DIN2_t(n6320_t),
    .Q(n4561),
    .Q_t(n4561_t)
  );


  nor2s3
  U3568
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4562),
    .DIN2_t(n4562_t),
    .Q(WX11660),
    .Q_t(WX11660_t)
  );


  xor2s3
  U3569
  (
    .DIN1(n6311),
    .DIN1_t(n6311_t),
    .DIN2(n6315),
    .DIN2_t(n6315_t),
    .Q(n4562),
    .Q_t(n4562_t)
  );


  nor2s3
  U3570
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4563),
    .DIN2_t(n4563_t),
    .Q(WX11658),
    .Q_t(WX11658_t)
  );


  xor2s3
  U3571
  (
    .DIN1(n6306),
    .DIN1_t(n6306_t),
    .DIN2(n6310),
    .DIN2_t(n6310_t),
    .Q(n4563),
    .Q_t(n4563_t)
  );


  nor2s3
  U3572
  (
    .DIN1(n6807),
    .DIN1_t(n6807_t),
    .DIN2(n4564),
    .DIN2_t(n4564_t),
    .Q(WX11656),
    .Q_t(WX11656_t)
  );


  xor2s3
  U3573
  (
    .DIN1(n6301),
    .DIN1_t(n6301_t),
    .DIN2(n6305),
    .DIN2_t(n6305_t),
    .Q(n4564),
    .Q_t(n4564_t)
  );


  nor2s3
  U3574
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4565),
    .DIN2_t(n4565_t),
    .Q(WX11654),
    .Q_t(WX11654_t)
  );


  xor2s3
  U3575
  (
    .DIN1(n6296),
    .DIN1_t(n6296_t),
    .DIN2(n6300),
    .DIN2_t(n6300_t),
    .Q(n4565),
    .Q_t(n4565_t)
  );


  nor2s3
  U3576
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4566),
    .DIN2_t(n4566_t),
    .Q(WX11652),
    .Q_t(WX11652_t)
  );


  xor2s3
  U3577
  (
    .DIN1(n6291),
    .DIN1_t(n6291_t),
    .DIN2(n6295),
    .DIN2_t(n6295_t),
    .Q(n4566),
    .Q_t(n4566_t)
  );


  nor2s3
  U3578
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4567),
    .DIN2_t(n4567_t),
    .Q(WX11650),
    .Q_t(WX11650_t)
  );


  xor2s3
  U3579
  (
    .DIN1(n6285),
    .DIN1_t(n6285_t),
    .DIN2(n6290),
    .DIN2_t(n6290_t),
    .Q(n4567),
    .Q_t(n4567_t)
  );


  nor2s3
  U3580
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4568),
    .DIN2_t(n4568_t),
    .Q(WX11648),
    .Q_t(WX11648_t)
  );


  xor2s3
  U3581
  (
    .DIN1(n6280),
    .DIN1_t(n6280_t),
    .DIN2(n6284),
    .DIN2_t(n6284_t),
    .Q(n4568),
    .Q_t(n4568_t)
  );


  nor2s3
  U3582
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4569),
    .DIN2_t(n4569_t),
    .Q(WX11646),
    .Q_t(WX11646_t)
  );


  xor2s3
  U3583
  (
    .DIN1(n6275),
    .DIN1_t(n6275_t),
    .DIN2(n6279),
    .DIN2_t(n6279_t),
    .Q(n4569),
    .Q_t(n4569_t)
  );


  nor2s3
  U3584
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4570),
    .DIN2_t(n4570_t),
    .Q(WX11644),
    .Q_t(WX11644_t)
  );


  xor2s3
  U3585
  (
    .DIN1(n6270),
    .DIN1_t(n6270_t),
    .DIN2(n6274),
    .DIN2_t(n6274_t),
    .Q(n4570),
    .Q_t(n4570_t)
  );


  nor2s3
  U3586
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4571),
    .DIN2_t(n4571_t),
    .Q(WX11642),
    .Q_t(WX11642_t)
  );


  xor2s3
  U3587
  (
    .DIN1(n6265),
    .DIN1_t(n6265_t),
    .DIN2(n6269),
    .DIN2_t(n6269_t),
    .Q(n4571),
    .Q_t(n4571_t)
  );


  nor2s3
  U3588
  (
    .DIN1(n4572),
    .DIN1_t(n4572_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX11640),
    .Q_t(WX11640_t)
  );


  xor2s3
  U3589
  (
    .DIN1(n1729),
    .DIN1_t(n1729_t),
    .DIN2(n4573),
    .DIN2_t(n4573_t),
    .Q(n4572),
    .Q_t(n4572_t)
  );


  xor2s3
  U3590
  (
    .DIN1(n6260),
    .DIN1_t(n6260_t),
    .DIN2(n6264),
    .DIN2_t(n6264_t),
    .Q(n4573),
    .Q_t(n4573_t)
  );


  nor2s3
  U3591
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4574),
    .DIN2_t(n4574_t),
    .Q(WX11638),
    .Q_t(WX11638_t)
  );


  xor2s3
  U3592
  (
    .DIN1(n6256),
    .DIN1_t(n6256_t),
    .DIN2(n3332),
    .DIN2_t(n3332_t),
    .Q(n4574),
    .Q_t(n4574_t)
  );


  nor2s3
  U3593
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4575),
    .DIN2_t(n4575_t),
    .Q(WX11636),
    .Q_t(WX11636_t)
  );


  xor2s3
  U3594
  (
    .DIN1(n6252),
    .DIN1_t(n6252_t),
    .DIN2(n3331),
    .DIN2_t(n3331_t),
    .Q(n4575),
    .Q_t(n4575_t)
  );


  nor2s3
  U3595
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4576),
    .DIN2_t(n4576_t),
    .Q(WX11634),
    .Q_t(WX11634_t)
  );


  xor2s3
  U3596
  (
    .DIN1(n6248),
    .DIN1_t(n6248_t),
    .DIN2(n3330),
    .DIN2_t(n3330_t),
    .Q(n4576),
    .Q_t(n4576_t)
  );


  nor2s3
  U3597
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4577),
    .DIN2_t(n4577_t),
    .Q(WX11632),
    .Q_t(WX11632_t)
  );


  xor2s3
  U3598
  (
    .DIN1(n6244),
    .DIN1_t(n6244_t),
    .DIN2(n3329),
    .DIN2_t(n3329_t),
    .Q(n4577),
    .Q_t(n4577_t)
  );


  nor2s3
  U3599
  (
    .DIN1(n4578),
    .DIN1_t(n4578_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX11630),
    .Q_t(WX11630_t)
  );


  xnr2s3
  U3600
  (
    .DIN1(n3328),
    .DIN1_t(n3328_t),
    .DIN2(n4579),
    .DIN2_t(n4579_t),
    .Q(n4578),
    .Q_t(n4578_t)
  );


  xor2s3
  U3601
  (
    .DIN1(n6240),
    .DIN1_t(n6240_t),
    .DIN2(n6337),
    .DIN2_t(n6337_t),
    .Q(n4579),
    .Q_t(n4579_t)
  );


  nor2s3
  U3602
  (
    .DIN1(n6808),
    .DIN1_t(n6808_t),
    .DIN2(n4580),
    .DIN2_t(n4580_t),
    .Q(WX11628),
    .Q_t(WX11628_t)
  );


  xor2s3
  U3603
  (
    .DIN1(n6236),
    .DIN1_t(n6236_t),
    .DIN2(n3327),
    .DIN2_t(n3327_t),
    .Q(n4580),
    .Q_t(n4580_t)
  );


  nor2s3
  U3604
  (
    .DIN1(n6788),
    .DIN1_t(n6788_t),
    .DIN2(n4581),
    .DIN2_t(n4581_t),
    .Q(WX11626),
    .Q_t(WX11626_t)
  );


  xor2s3
  U3605
  (
    .DIN1(n6232),
    .DIN1_t(n6232_t),
    .DIN2(n3326),
    .DIN2_t(n3326_t),
    .Q(n4581),
    .Q_t(n4581_t)
  );


  nor2s3
  U3606
  (
    .DIN1(n6788),
    .DIN1_t(n6788_t),
    .DIN2(n4582),
    .DIN2_t(n4582_t),
    .Q(WX11624),
    .Q_t(WX11624_t)
  );


  xor2s3
  U3607
  (
    .DIN1(n6228),
    .DIN1_t(n6228_t),
    .DIN2(n3325),
    .DIN2_t(n3325_t),
    .Q(n4582),
    .Q_t(n4582_t)
  );


  nor2s3
  U3608
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n4583),
    .DIN2_t(n4583_t),
    .Q(WX11622),
    .Q_t(WX11622_t)
  );


  xor2s3
  U3609
  (
    .DIN1(n6224),
    .DIN1_t(n6224_t),
    .DIN2(n3324),
    .DIN2_t(n3324_t),
    .Q(n4583),
    .Q_t(n4583_t)
  );


  nor2s3
  U3610
  (
    .DIN1(n6788),
    .DIN1_t(n6788_t),
    .DIN2(n4584),
    .DIN2_t(n4584_t),
    .Q(WX11620),
    .Q_t(WX11620_t)
  );


  xor2s3
  U3611
  (
    .DIN1(n6220),
    .DIN1_t(n6220_t),
    .DIN2(n3323),
    .DIN2_t(n3323_t),
    .Q(n4584),
    .Q_t(n4584_t)
  );


  nor2s3
  U3612
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n4585),
    .DIN2_t(n4585_t),
    .Q(WX11618),
    .Q_t(WX11618_t)
  );


  xor2s3
  U3613
  (
    .DIN1(n6216),
    .DIN1_t(n6216_t),
    .DIN2(n3322),
    .DIN2_t(n3322_t),
    .Q(n4585),
    .Q_t(n4585_t)
  );


  nor2s3
  U3614
  (
    .DIN1(n4586),
    .DIN1_t(n4586_t),
    .DIN2(n6776),
    .DIN2_t(n6776_t),
    .Q(WX11616),
    .Q_t(WX11616_t)
  );


  xnr2s3
  U3615
  (
    .DIN1(n3321),
    .DIN1_t(n3321_t),
    .DIN2(n4587),
    .DIN2_t(n4587_t),
    .Q(n4586),
    .Q_t(n4586_t)
  );


  xor2s3
  U3616
  (
    .DIN1(n6212),
    .DIN1_t(n6212_t),
    .DIN2(n6337),
    .DIN2_t(n6337_t),
    .Q(n4587),
    .Q_t(n4587_t)
  );


  nor2s3
  U3617
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n4588),
    .DIN2_t(n4588_t),
    .Q(WX11614),
    .Q_t(WX11614_t)
  );


  xor2s3
  U3618
  (
    .DIN1(n6208),
    .DIN1_t(n6208_t),
    .DIN2(n3320),
    .DIN2_t(n3320_t),
    .Q(n4588),
    .Q_t(n4588_t)
  );


  nor2s3
  U3619
  (
    .DIN1(n6788),
    .DIN1_t(n6788_t),
    .DIN2(n4589),
    .DIN2_t(n4589_t),
    .Q(WX11612),
    .Q_t(WX11612_t)
  );


  xor2s3
  U3620
  (
    .DIN1(n6204),
    .DIN1_t(n6204_t),
    .DIN2(n3319),
    .DIN2_t(n3319_t),
    .Q(n4589),
    .Q_t(n4589_t)
  );


  nor2s3
  U3621
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n4590),
    .DIN2_t(n4590_t),
    .Q(WX11610),
    .Q_t(WX11610_t)
  );


  xor2s3
  U3622
  (
    .DIN1(n6200),
    .DIN1_t(n6200_t),
    .DIN2(n3318),
    .DIN2_t(n3318_t),
    .Q(n4590),
    .Q_t(n4590_t)
  );


  nor2s3
  U3623
  (
    .DIN1(n6788),
    .DIN1_t(n6788_t),
    .DIN2(n4591),
    .DIN2_t(n4591_t),
    .Q(WX11608),
    .Q_t(WX11608_t)
  );


  xor2s3
  U3624
  (
    .DIN1(n6337),
    .DIN1_t(n6337_t),
    .DIN2(n3317),
    .DIN2_t(n3317_t),
    .Q(n4591),
    .Q_t(n4591_t)
  );


  nor2s3
  U3625
  (
    .DIN1(n6199),
    .DIN1_t(n6199_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX11242),
    .Q_t(WX11242_t)
  );


  nor2s3
  U3626
  (
    .DIN1(n6203),
    .DIN1_t(n6203_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX11240),
    .Q_t(WX11240_t)
  );


  nor2s3
  U3627
  (
    .DIN1(n6207),
    .DIN1_t(n6207_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX11238),
    .Q_t(WX11238_t)
  );


  nor2s3
  U3628
  (
    .DIN1(n6211),
    .DIN1_t(n6211_t),
    .DIN2(n6774),
    .DIN2_t(n6774_t),
    .Q(WX11236),
    .Q_t(WX11236_t)
  );


  nor2s3
  U3629
  (
    .DIN1(n6215),
    .DIN1_t(n6215_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11234),
    .Q_t(WX11234_t)
  );


  nor2s3
  U3630
  (
    .DIN1(n6219),
    .DIN1_t(n6219_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11232),
    .Q_t(WX11232_t)
  );


  nor2s3
  U3631
  (
    .DIN1(n6223),
    .DIN1_t(n6223_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11230),
    .Q_t(WX11230_t)
  );


  nor2s3
  U3632
  (
    .DIN1(n6227),
    .DIN1_t(n6227_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11228),
    .Q_t(WX11228_t)
  );


  nor2s3
  U3633
  (
    .DIN1(n6231),
    .DIN1_t(n6231_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11226),
    .Q_t(WX11226_t)
  );


  nor2s3
  U3634
  (
    .DIN1(n6235),
    .DIN1_t(n6235_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11224),
    .Q_t(WX11224_t)
  );


  nor2s3
  U3635
  (
    .DIN1(n6239),
    .DIN1_t(n6239_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11222),
    .Q_t(WX11222_t)
  );


  nor2s3
  U3636
  (
    .DIN1(n6243),
    .DIN1_t(n6243_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11220),
    .Q_t(WX11220_t)
  );


  nor2s3
  U3637
  (
    .DIN1(n6247),
    .DIN1_t(n6247_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11218),
    .Q_t(WX11218_t)
  );


  nor2s3
  U3638
  (
    .DIN1(n6251),
    .DIN1_t(n6251_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11216),
    .Q_t(WX11216_t)
  );


  nor2s3
  U3639
  (
    .DIN1(n6255),
    .DIN1_t(n6255_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11214),
    .Q_t(WX11214_t)
  );


  nor2s3
  U3640
  (
    .DIN1(n6259),
    .DIN1_t(n6259_t),
    .DIN2(n6773),
    .DIN2_t(n6773_t),
    .Q(WX11212),
    .Q_t(WX11212_t)
  );


  nor2s3
  U3641
  (
    .DIN1(n6263),
    .DIN1_t(n6263_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11210),
    .Q_t(WX11210_t)
  );


  nor2s3
  U3642
  (
    .DIN1(n6268),
    .DIN1_t(n6268_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11208),
    .Q_t(WX11208_t)
  );


  nor2s3
  U3643
  (
    .DIN1(n6273),
    .DIN1_t(n6273_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11206),
    .Q_t(WX11206_t)
  );


  nor2s3
  U3644
  (
    .DIN1(n6278),
    .DIN1_t(n6278_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11204),
    .Q_t(WX11204_t)
  );


  nor2s3
  U3645
  (
    .DIN1(n6283),
    .DIN1_t(n6283_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11202),
    .Q_t(WX11202_t)
  );


  nor2s3
  U3646
  (
    .DIN1(n6289),
    .DIN1_t(n6289_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11200),
    .Q_t(WX11200_t)
  );


  nor2s3
  U3647
  (
    .DIN1(n6294),
    .DIN1_t(n6294_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11198),
    .Q_t(WX11198_t)
  );


  nor2s3
  U3648
  (
    .DIN1(n6299),
    .DIN1_t(n6299_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11196),
    .Q_t(WX11196_t)
  );


  nor2s3
  U3649
  (
    .DIN1(n6304),
    .DIN1_t(n6304_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11194),
    .Q_t(WX11194_t)
  );


  nor2s3
  U3650
  (
    .DIN1(n6309),
    .DIN1_t(n6309_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11192),
    .Q_t(WX11192_t)
  );


  nor2s3
  U3651
  (
    .DIN1(n6314),
    .DIN1_t(n6314_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11190),
    .Q_t(WX11190_t)
  );


  nor2s3
  U3652
  (
    .DIN1(n6319),
    .DIN1_t(n6319_t),
    .DIN2(n6772),
    .DIN2_t(n6772_t),
    .Q(WX11188),
    .Q_t(WX11188_t)
  );


  nor2s3
  U3653
  (
    .DIN1(n6324),
    .DIN1_t(n6324_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX11186),
    .Q_t(WX11186_t)
  );


  nor2s3
  U3654
  (
    .DIN1(n6329),
    .DIN1_t(n6329_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX11184),
    .Q_t(WX11184_t)
  );


  nor2s3
  U3655
  (
    .DIN1(n6334),
    .DIN1_t(n6334_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX11182),
    .Q_t(WX11182_t)
  );


  nor2s3
  U3656
  (
    .DIN1(n6340),
    .DIN1_t(n6340_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX11180),
    .Q_t(WX11180_t)
  );


  and2s3
  U3657
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6198),
    .DIN2_t(n6198_t),
    .Q(WX11178),
    .Q_t(WX11178_t)
  );


  and2s3
  U3658
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6202),
    .DIN2_t(n6202_t),
    .Q(WX11176),
    .Q_t(WX11176_t)
  );


  and2s3
  U3659
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6206),
    .DIN2_t(n6206_t),
    .Q(WX11174),
    .Q_t(WX11174_t)
  );


  and2s3
  U3660
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6210),
    .DIN2_t(n6210_t),
    .Q(WX11172),
    .Q_t(WX11172_t)
  );


  and2s3
  U3661
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6214),
    .DIN2_t(n6214_t),
    .Q(WX11170),
    .Q_t(WX11170_t)
  );


  and2s3
  U3662
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6218),
    .DIN2_t(n6218_t),
    .Q(WX11168),
    .Q_t(WX11168_t)
  );


  and2s3
  U3663
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6222),
    .DIN2_t(n6222_t),
    .Q(WX11166),
    .Q_t(WX11166_t)
  );


  and2s3
  U3664
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6226),
    .DIN2_t(n6226_t),
    .Q(WX11164),
    .Q_t(WX11164_t)
  );


  and2s3
  U3665
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6230),
    .DIN2_t(n6230_t),
    .Q(WX11162),
    .Q_t(WX11162_t)
  );


  and2s3
  U3666
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6234),
    .DIN2_t(n6234_t),
    .Q(WX11160),
    .Q_t(WX11160_t)
  );


  and2s3
  U3667
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6238),
    .DIN2_t(n6238_t),
    .Q(WX11158),
    .Q_t(WX11158_t)
  );


  and2s3
  U3668
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6242),
    .DIN2_t(n6242_t),
    .Q(WX11156),
    .Q_t(WX11156_t)
  );


  and2s3
  U3669
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6246),
    .DIN2_t(n6246_t),
    .Q(WX11154),
    .Q_t(WX11154_t)
  );


  and2s3
  U3670
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6250),
    .DIN2_t(n6250_t),
    .Q(WX11152),
    .Q_t(WX11152_t)
  );


  and2s3
  U3671
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6254),
    .DIN2_t(n6254_t),
    .Q(WX11150),
    .Q_t(WX11150_t)
  );


  and2s3
  U3672
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6258),
    .DIN2_t(n6258_t),
    .Q(WX11148),
    .Q_t(WX11148_t)
  );


  and2s3
  U3673
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6262),
    .DIN2_t(n6262_t),
    .Q(WX11146),
    .Q_t(WX11146_t)
  );


  and2s3
  U3674
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6267),
    .DIN2_t(n6267_t),
    .Q(WX11144),
    .Q_t(WX11144_t)
  );


  and2s3
  U3675
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6272),
    .DIN2_t(n6272_t),
    .Q(WX11142),
    .Q_t(WX11142_t)
  );


  and2s3
  U3676
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6277),
    .DIN2_t(n6277_t),
    .Q(WX11140),
    .Q_t(WX11140_t)
  );


  and2s3
  U3677
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6282),
    .DIN2_t(n6282_t),
    .Q(WX11138),
    .Q_t(WX11138_t)
  );


  and2s3
  U3678
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6288),
    .DIN2_t(n6288_t),
    .Q(WX11136),
    .Q_t(WX11136_t)
  );


  and2s3
  U3679
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6293),
    .DIN2_t(n6293_t),
    .Q(WX11134),
    .Q_t(WX11134_t)
  );


  and2s3
  U3680
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6298),
    .DIN2_t(n6298_t),
    .Q(WX11132),
    .Q_t(WX11132_t)
  );


  and2s3
  U3681
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6303),
    .DIN2_t(n6303_t),
    .Q(WX11130),
    .Q_t(WX11130_t)
  );


  and2s3
  U3682
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6308),
    .DIN2_t(n6308_t),
    .Q(WX11128),
    .Q_t(WX11128_t)
  );


  and2s3
  U3683
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6313),
    .DIN2_t(n6313_t),
    .Q(WX11126),
    .Q_t(WX11126_t)
  );


  and2s3
  U3684
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6318),
    .DIN2_t(n6318_t),
    .Q(WX11124),
    .Q_t(WX11124_t)
  );


  and2s3
  U3685
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6323),
    .DIN2_t(n6323_t),
    .Q(WX11122),
    .Q_t(WX11122_t)
  );


  and2s3
  U3686
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6328),
    .DIN2_t(n6328_t),
    .Q(WX11120),
    .Q_t(WX11120_t)
  );


  and2s3
  U3687
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6333),
    .DIN2_t(n6333_t),
    .Q(WX11118),
    .Q_t(WX11118_t)
  );


  and2s3
  U3688
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6339),
    .DIN2_t(n6339_t),
    .Q(WX11116),
    .Q_t(WX11116_t)
  );


  nor2s3
  U3689
  (
    .DIN1(n6197),
    .DIN1_t(n6197_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX11114),
    .Q_t(WX11114_t)
  );


  nor2s3
  U3690
  (
    .DIN1(n6201),
    .DIN1_t(n6201_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX11112),
    .Q_t(WX11112_t)
  );


  nor2s3
  U3691
  (
    .DIN1(n6205),
    .DIN1_t(n6205_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX11110),
    .Q_t(WX11110_t)
  );


  nor2s3
  U3692
  (
    .DIN1(n6209),
    .DIN1_t(n6209_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX11108),
    .Q_t(WX11108_t)
  );


  nor2s3
  U3693
  (
    .DIN1(n6213),
    .DIN1_t(n6213_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX11106),
    .Q_t(WX11106_t)
  );


  nor2s3
  U3694
  (
    .DIN1(n6217),
    .DIN1_t(n6217_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX11104),
    .Q_t(WX11104_t)
  );


  nor2s3
  U3695
  (
    .DIN1(n6221),
    .DIN1_t(n6221_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX11102),
    .Q_t(WX11102_t)
  );


  nor2s3
  U3696
  (
    .DIN1(n6225),
    .DIN1_t(n6225_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11100),
    .Q_t(WX11100_t)
  );


  nor2s3
  U3697
  (
    .DIN1(n6229),
    .DIN1_t(n6229_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11098),
    .Q_t(WX11098_t)
  );


  nor2s3
  U3698
  (
    .DIN1(n6233),
    .DIN1_t(n6233_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11096),
    .Q_t(WX11096_t)
  );


  nor2s3
  U3699
  (
    .DIN1(n6237),
    .DIN1_t(n6237_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11094),
    .Q_t(WX11094_t)
  );


  nor2s3
  U3700
  (
    .DIN1(n6241),
    .DIN1_t(n6241_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11092),
    .Q_t(WX11092_t)
  );


  nor2s3
  U3701
  (
    .DIN1(n6245),
    .DIN1_t(n6245_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11090),
    .Q_t(WX11090_t)
  );


  nor2s3
  U3702
  (
    .DIN1(n6249),
    .DIN1_t(n6249_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11088),
    .Q_t(WX11088_t)
  );


  nor2s3
  U3703
  (
    .DIN1(n6253),
    .DIN1_t(n6253_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11086),
    .Q_t(WX11086_t)
  );


  nor2s3
  U3704
  (
    .DIN1(n6257),
    .DIN1_t(n6257_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11084),
    .Q_t(WX11084_t)
  );


  nor2s3
  U3705
  (
    .DIN1(n6261),
    .DIN1_t(n6261_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11082),
    .Q_t(WX11082_t)
  );


  nor2s3
  U3706
  (
    .DIN1(n6266),
    .DIN1_t(n6266_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11080),
    .Q_t(WX11080_t)
  );


  nor2s3
  U3707
  (
    .DIN1(n6271),
    .DIN1_t(n6271_t),
    .DIN2(n6770),
    .DIN2_t(n6770_t),
    .Q(WX11078),
    .Q_t(WX11078_t)
  );


  nor2s3
  U3708
  (
    .DIN1(n6276),
    .DIN1_t(n6276_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11076),
    .Q_t(WX11076_t)
  );


  nor2s3
  U3709
  (
    .DIN1(n6281),
    .DIN1_t(n6281_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11074),
    .Q_t(WX11074_t)
  );


  nor2s3
  U3710
  (
    .DIN1(n6287),
    .DIN1_t(n6287_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11072),
    .Q_t(WX11072_t)
  );


  nor2s3
  U3711
  (
    .DIN1(n6292),
    .DIN1_t(n6292_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11070),
    .Q_t(WX11070_t)
  );


  nor2s3
  U3712
  (
    .DIN1(n6297),
    .DIN1_t(n6297_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11068),
    .Q_t(WX11068_t)
  );


  nor2s3
  U3713
  (
    .DIN1(n6302),
    .DIN1_t(n6302_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11066),
    .Q_t(WX11066_t)
  );


  nor2s3
  U3714
  (
    .DIN1(n6307),
    .DIN1_t(n6307_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11064),
    .Q_t(WX11064_t)
  );


  nor2s3
  U3715
  (
    .DIN1(n6312),
    .DIN1_t(n6312_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11062),
    .Q_t(WX11062_t)
  );


  nor2s3
  U3716
  (
    .DIN1(n6317),
    .DIN1_t(n6317_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11060),
    .Q_t(WX11060_t)
  );


  nor2s3
  U3717
  (
    .DIN1(n6322),
    .DIN1_t(n6322_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11058),
    .Q_t(WX11058_t)
  );


  nor2s3
  U3718
  (
    .DIN1(n6327),
    .DIN1_t(n6327_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11056),
    .Q_t(WX11056_t)
  );


  nor2s3
  U3719
  (
    .DIN1(n6332),
    .DIN1_t(n6332_t),
    .DIN2(n6769),
    .DIN2_t(n6769_t),
    .Q(WX11054),
    .Q_t(WX11054_t)
  );


  nor2s3
  U3720
  (
    .DIN1(n6338),
    .DIN1_t(n6338_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX11052),
    .Q_t(WX11052_t)
  );


  nnd4s2
  U3721
  (
    .DIN1(n4592),
    .DIN1_t(n4592_t),
    .DIN2(n4593),
    .DIN2_t(n4593_t),
    .DIN3(n4594),
    .DIN3_t(n4594_t),
    .DIN4(n4595),
    .DIN4_t(n4595_t),
    .Q(WX11050),
    .Q_t(WX11050_t)
  );


  nnd2s3
  U3722
  (
    .DIN1(n2315),
    .DIN1_t(n2315_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4595),
    .Q_t(n4595_t)
  );


  xor2s3
  U3723
  (
    .DIN1(n4596),
    .DIN1_t(n4596_t),
    .DIN2(n4597),
    .DIN2_t(n4597_t),
    .Q(n2315),
    .Q_t(n2315_t)
  );


  xor2s3
  U3724
  (
    .DIN1(n6197),
    .DIN1_t(n6197_t),
    .DIN2(n6198),
    .DIN2_t(n6198_t),
    .Q(n4597),
    .Q_t(n4597_t)
  );


  xnr2s3
  U3725
  (
    .DIN1(n3317),
    .DIN1_t(n3317_t),
    .DIN2(n6199),
    .DIN2_t(n6199_t),
    .Q(n4596),
    .Q_t(n4596_t)
  );


  nnd2s3
  U3726
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n1761),
    .DIN2_t(n1761_t),
    .Q(n4594),
    .Q_t(n4594_t)
  );


  nnd2s3
  U3727
  (
    .DIN1(DATA_0_0),
    .DIN1_t(DATA_0_0_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4593),
    .Q_t(n4593_t)
  );


  nnd2s3
  U3728
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n1760),
    .DIN2_t(n1760_t),
    .Q(n4592),
    .Q_t(n4592_t)
  );


  nnd4s2
  U3729
  (
    .DIN1(n4598),
    .DIN1_t(n4598_t),
    .DIN2(n4599),
    .DIN2_t(n4599_t),
    .DIN3(n4600),
    .DIN3_t(n4600_t),
    .DIN4(n4601),
    .DIN4_t(n4601_t),
    .Q(WX11048),
    .Q_t(WX11048_t)
  );


  nnd2s3
  U3730
  (
    .DIN1(n2323),
    .DIN1_t(n2323_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4601),
    .Q_t(n4601_t)
  );


  xor2s3
  U3731
  (
    .DIN1(n4602),
    .DIN1_t(n4602_t),
    .DIN2(n4603),
    .DIN2_t(n4603_t),
    .Q(n2323),
    .Q_t(n2323_t)
  );


  xor2s3
  U3732
  (
    .DIN1(n6201),
    .DIN1_t(n6201_t),
    .DIN2(n6202),
    .DIN2_t(n6202_t),
    .Q(n4603),
    .Q_t(n4603_t)
  );


  xnr2s3
  U3733
  (
    .DIN1(n3318),
    .DIN1_t(n3318_t),
    .DIN2(n6203),
    .DIN2_t(n6203_t),
    .Q(n4602),
    .Q_t(n4602_t)
  );


  nnd2s3
  U3734
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n1762),
    .DIN2_t(n1762_t),
    .Q(n4600),
    .Q_t(n4600_t)
  );


  nnd2s3
  U3735
  (
    .DIN1(DATA_0_1),
    .DIN1_t(DATA_0_1_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4599),
    .Q_t(n4599_t)
  );


  nnd2s3
  U3736
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n1759),
    .DIN2_t(n1759_t),
    .Q(n4598),
    .Q_t(n4598_t)
  );


  nnd4s2
  U3737
  (
    .DIN1(n4604),
    .DIN1_t(n4604_t),
    .DIN2(n4605),
    .DIN2_t(n4605_t),
    .DIN3(n4606),
    .DIN3_t(n4606_t),
    .DIN4(n4607),
    .DIN4_t(n4607_t),
    .Q(WX11046),
    .Q_t(WX11046_t)
  );


  nnd2s3
  U3738
  (
    .DIN1(n2329),
    .DIN1_t(n2329_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4607),
    .Q_t(n4607_t)
  );


  xor2s3
  U3739
  (
    .DIN1(n4608),
    .DIN1_t(n4608_t),
    .DIN2(n4609),
    .DIN2_t(n4609_t),
    .Q(n2329),
    .Q_t(n2329_t)
  );


  xor2s3
  U3740
  (
    .DIN1(n6205),
    .DIN1_t(n6205_t),
    .DIN2(n6206),
    .DIN2_t(n6206_t),
    .Q(n4609),
    .Q_t(n4609_t)
  );


  xnr2s3
  U3741
  (
    .DIN1(n3319),
    .DIN1_t(n3319_t),
    .DIN2(n6207),
    .DIN2_t(n6207_t),
    .Q(n4608),
    .Q_t(n4608_t)
  );


  nnd2s3
  U3742
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n1763),
    .DIN2_t(n1763_t),
    .Q(n4606),
    .Q_t(n4606_t)
  );


  nnd2s3
  U3743
  (
    .DIN1(DATA_0_2),
    .DIN1_t(DATA_0_2_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4605),
    .Q_t(n4605_t)
  );


  nnd2s3
  U3744
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n1758),
    .DIN2_t(n1758_t),
    .Q(n4604),
    .Q_t(n4604_t)
  );


  nnd4s2
  U3745
  (
    .DIN1(n4610),
    .DIN1_t(n4610_t),
    .DIN2(n4611),
    .DIN2_t(n4611_t),
    .DIN3(n4612),
    .DIN3_t(n4612_t),
    .DIN4(n4613),
    .DIN4_t(n4613_t),
    .Q(WX11044),
    .Q_t(WX11044_t)
  );


  nnd2s3
  U3746
  (
    .DIN1(n2335),
    .DIN1_t(n2335_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4613),
    .Q_t(n4613_t)
  );


  xor2s3
  U3747
  (
    .DIN1(n4614),
    .DIN1_t(n4614_t),
    .DIN2(n4615),
    .DIN2_t(n4615_t),
    .Q(n2335),
    .Q_t(n2335_t)
  );


  xor2s3
  U3748
  (
    .DIN1(n6209),
    .DIN1_t(n6209_t),
    .DIN2(n6210),
    .DIN2_t(n6210_t),
    .Q(n4615),
    .Q_t(n4615_t)
  );


  xnr2s3
  U3749
  (
    .DIN1(n3320),
    .DIN1_t(n3320_t),
    .DIN2(n6211),
    .DIN2_t(n6211_t),
    .Q(n4614),
    .Q_t(n4614_t)
  );


  nnd2s3
  U3750
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n1764),
    .DIN2_t(n1764_t),
    .Q(n4612),
    .Q_t(n4612_t)
  );


  nnd2s3
  U3751
  (
    .DIN1(DATA_0_3),
    .DIN1_t(DATA_0_3_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4611),
    .Q_t(n4611_t)
  );


  nnd2s3
  U3752
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n1757),
    .DIN2_t(n1757_t),
    .Q(n4610),
    .Q_t(n4610_t)
  );


  nnd4s2
  U3753
  (
    .DIN1(n4616),
    .DIN1_t(n4616_t),
    .DIN2(n4617),
    .DIN2_t(n4617_t),
    .DIN3(n4618),
    .DIN3_t(n4618_t),
    .DIN4(n4619),
    .DIN4_t(n4619_t),
    .Q(WX11042),
    .Q_t(WX11042_t)
  );


  nnd2s3
  U3754
  (
    .DIN1(n2341),
    .DIN1_t(n2341_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4619),
    .Q_t(n4619_t)
  );


  xor2s3
  U3755
  (
    .DIN1(n4620),
    .DIN1_t(n4620_t),
    .DIN2(n4621),
    .DIN2_t(n4621_t),
    .Q(n2341),
    .Q_t(n2341_t)
  );


  xor2s3
  U3756
  (
    .DIN1(n6213),
    .DIN1_t(n6213_t),
    .DIN2(n6214),
    .DIN2_t(n6214_t),
    .Q(n4621),
    .Q_t(n4621_t)
  );


  xnr2s3
  U3757
  (
    .DIN1(n3321),
    .DIN1_t(n3321_t),
    .DIN2(n6215),
    .DIN2_t(n6215_t),
    .Q(n4620),
    .Q_t(n4620_t)
  );


  nnd2s3
  U3758
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n1765),
    .DIN2_t(n1765_t),
    .Q(n4618),
    .Q_t(n4618_t)
  );


  nnd2s3
  U3759
  (
    .DIN1(DATA_0_4),
    .DIN1_t(DATA_0_4_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4617),
    .Q_t(n4617_t)
  );


  nnd2s3
  U3760
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n1756),
    .DIN2_t(n1756_t),
    .Q(n4616),
    .Q_t(n4616_t)
  );


  nnd4s2
  U3761
  (
    .DIN1(n4622),
    .DIN1_t(n4622_t),
    .DIN2(n4623),
    .DIN2_t(n4623_t),
    .DIN3(n4624),
    .DIN3_t(n4624_t),
    .DIN4(n4625),
    .DIN4_t(n4625_t),
    .Q(WX11040),
    .Q_t(WX11040_t)
  );


  nnd2s3
  U3762
  (
    .DIN1(n2347),
    .DIN1_t(n2347_t),
    .DIN2(n6669),
    .DIN2_t(n6669_t),
    .Q(n4625),
    .Q_t(n4625_t)
  );


  xor2s3
  U3763
  (
    .DIN1(n4626),
    .DIN1_t(n4626_t),
    .DIN2(n4627),
    .DIN2_t(n4627_t),
    .Q(n2347),
    .Q_t(n2347_t)
  );


  xor2s3
  U3764
  (
    .DIN1(n6217),
    .DIN1_t(n6217_t),
    .DIN2(n6218),
    .DIN2_t(n6218_t),
    .Q(n4627),
    .Q_t(n4627_t)
  );


  xnr2s3
  U3765
  (
    .DIN1(n3322),
    .DIN1_t(n3322_t),
    .DIN2(n6219),
    .DIN2_t(n6219_t),
    .Q(n4626),
    .Q_t(n4626_t)
  );


  nnd2s3
  U3766
  (
    .DIN1(n6596),
    .DIN1_t(n6596_t),
    .DIN2(n1766),
    .DIN2_t(n1766_t),
    .Q(n4624),
    .Q_t(n4624_t)
  );


  nnd2s3
  U3767
  (
    .DIN1(DATA_0_5),
    .DIN1_t(DATA_0_5_t),
    .DIN2(n6638),
    .DIN2_t(n6638_t),
    .Q(n4623),
    .Q_t(n4623_t)
  );


  nnd2s3
  U3768
  (
    .DIN1(n6565),
    .DIN1_t(n6565_t),
    .DIN2(n1755),
    .DIN2_t(n1755_t),
    .Q(n4622),
    .Q_t(n4622_t)
  );


  nnd4s2
  U3769
  (
    .DIN1(n4628),
    .DIN1_t(n4628_t),
    .DIN2(n4629),
    .DIN2_t(n4629_t),
    .DIN3(n4630),
    .DIN3_t(n4630_t),
    .DIN4(n4631),
    .DIN4_t(n4631_t),
    .Q(WX11038),
    .Q_t(WX11038_t)
  );


  nnd2s3
  U3770
  (
    .DIN1(n2353),
    .DIN1_t(n2353_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4631),
    .Q_t(n4631_t)
  );


  xor2s3
  U3771
  (
    .DIN1(n4632),
    .DIN1_t(n4632_t),
    .DIN2(n4633),
    .DIN2_t(n4633_t),
    .Q(n2353),
    .Q_t(n2353_t)
  );


  xor2s3
  U3772
  (
    .DIN1(n6221),
    .DIN1_t(n6221_t),
    .DIN2(n6222),
    .DIN2_t(n6222_t),
    .Q(n4633),
    .Q_t(n4633_t)
  );


  xnr2s3
  U3773
  (
    .DIN1(n3323),
    .DIN1_t(n3323_t),
    .DIN2(n6223),
    .DIN2_t(n6223_t),
    .Q(n4632),
    .Q_t(n4632_t)
  );


  nnd2s3
  U3774
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1767),
    .DIN2_t(n1767_t),
    .Q(n4630),
    .Q_t(n4630_t)
  );


  nnd2s3
  U3775
  (
    .DIN1(DATA_0_6),
    .DIN1_t(DATA_0_6_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4629),
    .Q_t(n4629_t)
  );


  nnd2s3
  U3776
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1754),
    .DIN2_t(n1754_t),
    .Q(n4628),
    .Q_t(n4628_t)
  );


  nnd4s2
  U3777
  (
    .DIN1(n4634),
    .DIN1_t(n4634_t),
    .DIN2(n4635),
    .DIN2_t(n4635_t),
    .DIN3(n4636),
    .DIN3_t(n4636_t),
    .DIN4(n4637),
    .DIN4_t(n4637_t),
    .Q(WX11036),
    .Q_t(WX11036_t)
  );


  nnd2s3
  U3778
  (
    .DIN1(n2359),
    .DIN1_t(n2359_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4637),
    .Q_t(n4637_t)
  );


  xor2s3
  U3779
  (
    .DIN1(n4638),
    .DIN1_t(n4638_t),
    .DIN2(n4639),
    .DIN2_t(n4639_t),
    .Q(n2359),
    .Q_t(n2359_t)
  );


  xor2s3
  U3780
  (
    .DIN1(n6225),
    .DIN1_t(n6225_t),
    .DIN2(n6226),
    .DIN2_t(n6226_t),
    .Q(n4639),
    .Q_t(n4639_t)
  );


  xnr2s3
  U3781
  (
    .DIN1(n3324),
    .DIN1_t(n3324_t),
    .DIN2(n6227),
    .DIN2_t(n6227_t),
    .Q(n4638),
    .Q_t(n4638_t)
  );


  nnd2s3
  U3782
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1768),
    .DIN2_t(n1768_t),
    .Q(n4636),
    .Q_t(n4636_t)
  );


  nnd2s3
  U3783
  (
    .DIN1(DATA_0_7),
    .DIN1_t(DATA_0_7_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4635),
    .Q_t(n4635_t)
  );


  nnd2s3
  U3784
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1753),
    .DIN2_t(n1753_t),
    .Q(n4634),
    .Q_t(n4634_t)
  );


  nnd4s2
  U3785
  (
    .DIN1(n4640),
    .DIN1_t(n4640_t),
    .DIN2(n4641),
    .DIN2_t(n4641_t),
    .DIN3(n4642),
    .DIN3_t(n4642_t),
    .DIN4(n4643),
    .DIN4_t(n4643_t),
    .Q(WX11034),
    .Q_t(WX11034_t)
  );


  nnd2s3
  U3786
  (
    .DIN1(n2365),
    .DIN1_t(n2365_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4643),
    .Q_t(n4643_t)
  );


  xor2s3
  U3787
  (
    .DIN1(n4644),
    .DIN1_t(n4644_t),
    .DIN2(n4645),
    .DIN2_t(n4645_t),
    .Q(n2365),
    .Q_t(n2365_t)
  );


  xor2s3
  U3788
  (
    .DIN1(n6229),
    .DIN1_t(n6229_t),
    .DIN2(n6230),
    .DIN2_t(n6230_t),
    .Q(n4645),
    .Q_t(n4645_t)
  );


  xnr2s3
  U3789
  (
    .DIN1(n3325),
    .DIN1_t(n3325_t),
    .DIN2(n6231),
    .DIN2_t(n6231_t),
    .Q(n4644),
    .Q_t(n4644_t)
  );


  nnd2s3
  U3790
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1769),
    .DIN2_t(n1769_t),
    .Q(n4642),
    .Q_t(n4642_t)
  );


  nnd2s3
  U3791
  (
    .DIN1(DATA_0_8),
    .DIN1_t(DATA_0_8_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4641),
    .Q_t(n4641_t)
  );


  nnd2s3
  U3792
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1752),
    .DIN2_t(n1752_t),
    .Q(n4640),
    .Q_t(n4640_t)
  );


  nnd4s2
  U3793
  (
    .DIN1(n4646),
    .DIN1_t(n4646_t),
    .DIN2(n4647),
    .DIN2_t(n4647_t),
    .DIN3(n4648),
    .DIN3_t(n4648_t),
    .DIN4(n4649),
    .DIN4_t(n4649_t),
    .Q(WX11032),
    .Q_t(WX11032_t)
  );


  nnd2s3
  U3794
  (
    .DIN1(n2371),
    .DIN1_t(n2371_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4649),
    .Q_t(n4649_t)
  );


  xor2s3
  U3795
  (
    .DIN1(n4650),
    .DIN1_t(n4650_t),
    .DIN2(n4651),
    .DIN2_t(n4651_t),
    .Q(n2371),
    .Q_t(n2371_t)
  );


  xor2s3
  U3796
  (
    .DIN1(n6233),
    .DIN1_t(n6233_t),
    .DIN2(n6234),
    .DIN2_t(n6234_t),
    .Q(n4651),
    .Q_t(n4651_t)
  );


  xnr2s3
  U3797
  (
    .DIN1(n3326),
    .DIN1_t(n3326_t),
    .DIN2(n6235),
    .DIN2_t(n6235_t),
    .Q(n4650),
    .Q_t(n4650_t)
  );


  nnd2s3
  U3798
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1770),
    .DIN2_t(n1770_t),
    .Q(n4648),
    .Q_t(n4648_t)
  );


  nnd2s3
  U3799
  (
    .DIN1(DATA_0_9),
    .DIN1_t(DATA_0_9_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4647),
    .Q_t(n4647_t)
  );


  nnd2s3
  U3800
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1751),
    .DIN2_t(n1751_t),
    .Q(n4646),
    .Q_t(n4646_t)
  );


  nnd4s2
  U3801
  (
    .DIN1(n4652),
    .DIN1_t(n4652_t),
    .DIN2(n4653),
    .DIN2_t(n4653_t),
    .DIN3(n4654),
    .DIN3_t(n4654_t),
    .DIN4(n4655),
    .DIN4_t(n4655_t),
    .Q(WX11030),
    .Q_t(WX11030_t)
  );


  nnd2s3
  U3802
  (
    .DIN1(n2377),
    .DIN1_t(n2377_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4655),
    .Q_t(n4655_t)
  );


  xor2s3
  U3803
  (
    .DIN1(n4656),
    .DIN1_t(n4656_t),
    .DIN2(n4657),
    .DIN2_t(n4657_t),
    .Q(n2377),
    .Q_t(n2377_t)
  );


  xor2s3
  U3804
  (
    .DIN1(n6237),
    .DIN1_t(n6237_t),
    .DIN2(n6238),
    .DIN2_t(n6238_t),
    .Q(n4657),
    .Q_t(n4657_t)
  );


  xnr2s3
  U3805
  (
    .DIN1(n3327),
    .DIN1_t(n3327_t),
    .DIN2(n6239),
    .DIN2_t(n6239_t),
    .Q(n4656),
    .Q_t(n4656_t)
  );


  nnd2s3
  U3806
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1771),
    .DIN2_t(n1771_t),
    .Q(n4654),
    .Q_t(n4654_t)
  );


  nnd2s3
  U3807
  (
    .DIN1(DATA_0_10),
    .DIN1_t(DATA_0_10_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4653),
    .Q_t(n4653_t)
  );


  nnd2s3
  U3808
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1750),
    .DIN2_t(n1750_t),
    .Q(n4652),
    .Q_t(n4652_t)
  );


  nnd4s2
  U3809
  (
    .DIN1(n4658),
    .DIN1_t(n4658_t),
    .DIN2(n4659),
    .DIN2_t(n4659_t),
    .DIN3(n4660),
    .DIN3_t(n4660_t),
    .DIN4(n4661),
    .DIN4_t(n4661_t),
    .Q(WX11028),
    .Q_t(WX11028_t)
  );


  nnd2s3
  U3810
  (
    .DIN1(n2383),
    .DIN1_t(n2383_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4661),
    .Q_t(n4661_t)
  );


  xor2s3
  U3811
  (
    .DIN1(n4662),
    .DIN1_t(n4662_t),
    .DIN2(n4663),
    .DIN2_t(n4663_t),
    .Q(n2383),
    .Q_t(n2383_t)
  );


  xor2s3
  U3812
  (
    .DIN1(n6241),
    .DIN1_t(n6241_t),
    .DIN2(n6242),
    .DIN2_t(n6242_t),
    .Q(n4663),
    .Q_t(n4663_t)
  );


  xnr2s3
  U3813
  (
    .DIN1(n3328),
    .DIN1_t(n3328_t),
    .DIN2(n6243),
    .DIN2_t(n6243_t),
    .Q(n4662),
    .Q_t(n4662_t)
  );


  nnd2s3
  U3814
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1772),
    .DIN2_t(n1772_t),
    .Q(n4660),
    .Q_t(n4660_t)
  );


  nnd2s3
  U3815
  (
    .DIN1(DATA_0_11),
    .DIN1_t(DATA_0_11_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4659),
    .Q_t(n4659_t)
  );


  nnd2s3
  U3816
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1749),
    .DIN2_t(n1749_t),
    .Q(n4658),
    .Q_t(n4658_t)
  );


  nnd4s2
  U3817
  (
    .DIN1(n4664),
    .DIN1_t(n4664_t),
    .DIN2(n4665),
    .DIN2_t(n4665_t),
    .DIN3(n4666),
    .DIN3_t(n4666_t),
    .DIN4(n4667),
    .DIN4_t(n4667_t),
    .Q(WX11026),
    .Q_t(WX11026_t)
  );


  nnd2s3
  U3818
  (
    .DIN1(n2389),
    .DIN1_t(n2389_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4667),
    .Q_t(n4667_t)
  );


  xor2s3
  U3819
  (
    .DIN1(n4668),
    .DIN1_t(n4668_t),
    .DIN2(n4669),
    .DIN2_t(n4669_t),
    .Q(n2389),
    .Q_t(n2389_t)
  );


  xor2s3
  U3820
  (
    .DIN1(n6245),
    .DIN1_t(n6245_t),
    .DIN2(n6246),
    .DIN2_t(n6246_t),
    .Q(n4669),
    .Q_t(n4669_t)
  );


  xnr2s3
  U3821
  (
    .DIN1(n3329),
    .DIN1_t(n3329_t),
    .DIN2(n6247),
    .DIN2_t(n6247_t),
    .Q(n4668),
    .Q_t(n4668_t)
  );


  nnd2s3
  U3822
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1773),
    .DIN2_t(n1773_t),
    .Q(n4666),
    .Q_t(n4666_t)
  );


  nnd2s3
  U3823
  (
    .DIN1(DATA_0_12),
    .DIN1_t(DATA_0_12_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4665),
    .Q_t(n4665_t)
  );


  nnd2s3
  U3824
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1748),
    .DIN2_t(n1748_t),
    .Q(n4664),
    .Q_t(n4664_t)
  );


  nnd4s2
  U3825
  (
    .DIN1(n4670),
    .DIN1_t(n4670_t),
    .DIN2(n4671),
    .DIN2_t(n4671_t),
    .DIN3(n4672),
    .DIN3_t(n4672_t),
    .DIN4(n4673),
    .DIN4_t(n4673_t),
    .Q(WX11024),
    .Q_t(WX11024_t)
  );


  nnd2s3
  U3826
  (
    .DIN1(n2395),
    .DIN1_t(n2395_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4673),
    .Q_t(n4673_t)
  );


  xor2s3
  U3827
  (
    .DIN1(n4674),
    .DIN1_t(n4674_t),
    .DIN2(n4675),
    .DIN2_t(n4675_t),
    .Q(n2395),
    .Q_t(n2395_t)
  );


  xor2s3
  U3828
  (
    .DIN1(n6249),
    .DIN1_t(n6249_t),
    .DIN2(n6250),
    .DIN2_t(n6250_t),
    .Q(n4675),
    .Q_t(n4675_t)
  );


  xnr2s3
  U3829
  (
    .DIN1(n3330),
    .DIN1_t(n3330_t),
    .DIN2(n6251),
    .DIN2_t(n6251_t),
    .Q(n4674),
    .Q_t(n4674_t)
  );


  nnd2s3
  U3830
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1774),
    .DIN2_t(n1774_t),
    .Q(n4672),
    .Q_t(n4672_t)
  );


  nnd2s3
  U3831
  (
    .DIN1(DATA_0_13),
    .DIN1_t(DATA_0_13_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4671),
    .Q_t(n4671_t)
  );


  nnd2s3
  U3832
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1747),
    .DIN2_t(n1747_t),
    .Q(n4670),
    .Q_t(n4670_t)
  );


  nnd4s2
  U3833
  (
    .DIN1(n4676),
    .DIN1_t(n4676_t),
    .DIN2(n4677),
    .DIN2_t(n4677_t),
    .DIN3(n4678),
    .DIN3_t(n4678_t),
    .DIN4(n4679),
    .DIN4_t(n4679_t),
    .Q(WX11022),
    .Q_t(WX11022_t)
  );


  nnd2s3
  U3834
  (
    .DIN1(n2401),
    .DIN1_t(n2401_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4679),
    .Q_t(n4679_t)
  );


  xor2s3
  U3835
  (
    .DIN1(n4680),
    .DIN1_t(n4680_t),
    .DIN2(n4681),
    .DIN2_t(n4681_t),
    .Q(n2401),
    .Q_t(n2401_t)
  );


  xor2s3
  U3836
  (
    .DIN1(n6253),
    .DIN1_t(n6253_t),
    .DIN2(n6254),
    .DIN2_t(n6254_t),
    .Q(n4681),
    .Q_t(n4681_t)
  );


  xnr2s3
  U3837
  (
    .DIN1(n3331),
    .DIN1_t(n3331_t),
    .DIN2(n6255),
    .DIN2_t(n6255_t),
    .Q(n4680),
    .Q_t(n4680_t)
  );


  nnd2s3
  U3838
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1775),
    .DIN2_t(n1775_t),
    .Q(n4678),
    .Q_t(n4678_t)
  );


  nnd2s3
  U3839
  (
    .DIN1(DATA_0_14),
    .DIN1_t(DATA_0_14_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4677),
    .Q_t(n4677_t)
  );


  nnd2s3
  U3840
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1746),
    .DIN2_t(n1746_t),
    .Q(n4676),
    .Q_t(n4676_t)
  );


  nnd4s2
  U3841
  (
    .DIN1(n4682),
    .DIN1_t(n4682_t),
    .DIN2(n4683),
    .DIN2_t(n4683_t),
    .DIN3(n4684),
    .DIN3_t(n4684_t),
    .DIN4(n4685),
    .DIN4_t(n4685_t),
    .Q(WX11020),
    .Q_t(WX11020_t)
  );


  nnd2s3
  U3842
  (
    .DIN1(n2407),
    .DIN1_t(n2407_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4685),
    .Q_t(n4685_t)
  );


  xor2s3
  U3843
  (
    .DIN1(n4686),
    .DIN1_t(n4686_t),
    .DIN2(n4687),
    .DIN2_t(n4687_t),
    .Q(n2407),
    .Q_t(n2407_t)
  );


  xor2s3
  U3844
  (
    .DIN1(n6257),
    .DIN1_t(n6257_t),
    .DIN2(n6258),
    .DIN2_t(n6258_t),
    .Q(n4687),
    .Q_t(n4687_t)
  );


  xnr2s3
  U3845
  (
    .DIN1(n3332),
    .DIN1_t(n3332_t),
    .DIN2(n6259),
    .DIN2_t(n6259_t),
    .Q(n4686),
    .Q_t(n4686_t)
  );


  nnd2s3
  U3846
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1776),
    .DIN2_t(n1776_t),
    .Q(n4684),
    .Q_t(n4684_t)
  );


  nnd2s3
  U3847
  (
    .DIN1(DATA_0_15),
    .DIN1_t(DATA_0_15_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4683),
    .Q_t(n4683_t)
  );


  nnd2s3
  U3848
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1745),
    .DIN2_t(n1745_t),
    .Q(n4682),
    .Q_t(n4682_t)
  );


  nnd4s2
  U3849
  (
    .DIN1(n4688),
    .DIN1_t(n4688_t),
    .DIN2(n4689),
    .DIN2_t(n4689_t),
    .DIN3(n4690),
    .DIN3_t(n4690_t),
    .DIN4(n4691),
    .DIN4_t(n4691_t),
    .Q(WX11018),
    .Q_t(WX11018_t)
  );


  nnd2s3
  U3850
  (
    .DIN1(n2413),
    .DIN1_t(n2413_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4691),
    .Q_t(n4691_t)
  );


  xor2s3
  U3851
  (
    .DIN1(n4692),
    .DIN1_t(n4692_t),
    .DIN2(n4693),
    .DIN2_t(n4693_t),
    .Q(n2413),
    .Q_t(n2413_t)
  );


  xor2s3
  U3852
  (
    .DIN1(n6263),
    .DIN1_t(n6263_t),
    .DIN2(n4694),
    .DIN2_t(n4694_t),
    .Q(n4693),
    .Q_t(n4693_t)
  );


  xor2s3
  U3853
  (
    .DIN1(n6261),
    .DIN1_t(n6261_t),
    .DIN2(n6262),
    .DIN2_t(n6262_t),
    .Q(n4694),
    .Q_t(n4694_t)
  );


  xor2s3
  U3854
  (
    .DIN1(n6264),
    .DIN1_t(n6264_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4692),
    .Q_t(n4692_t)
  );


  nnd2s3
  U3855
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1777),
    .DIN2_t(n1777_t),
    .Q(n4690),
    .Q_t(n4690_t)
  );


  nnd2s3
  U3856
  (
    .DIN1(DATA_0_16),
    .DIN1_t(DATA_0_16_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4689),
    .Q_t(n4689_t)
  );


  nnd2s3
  U3857
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1744),
    .DIN2_t(n1744_t),
    .Q(n4688),
    .Q_t(n4688_t)
  );


  nnd4s2
  U3858
  (
    .DIN1(n4695),
    .DIN1_t(n4695_t),
    .DIN2(n4696),
    .DIN2_t(n4696_t),
    .DIN3(n4697),
    .DIN3_t(n4697_t),
    .DIN4(n4698),
    .DIN4_t(n4698_t),
    .Q(WX11016),
    .Q_t(WX11016_t)
  );


  nnd2s3
  U3859
  (
    .DIN1(n2419),
    .DIN1_t(n2419_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4698),
    .Q_t(n4698_t)
  );


  xor2s3
  U3860
  (
    .DIN1(n4699),
    .DIN1_t(n4699_t),
    .DIN2(n4700),
    .DIN2_t(n4700_t),
    .Q(n2419),
    .Q_t(n2419_t)
  );


  xor2s3
  U3861
  (
    .DIN1(n6268),
    .DIN1_t(n6268_t),
    .DIN2(n4701),
    .DIN2_t(n4701_t),
    .Q(n4700),
    .Q_t(n4700_t)
  );


  xor2s3
  U3862
  (
    .DIN1(n6266),
    .DIN1_t(n6266_t),
    .DIN2(n6267),
    .DIN2_t(n6267_t),
    .Q(n4701),
    .Q_t(n4701_t)
  );


  xor2s3
  U3863
  (
    .DIN1(n6269),
    .DIN1_t(n6269_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4699),
    .Q_t(n4699_t)
  );


  nnd2s3
  U3864
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1778),
    .DIN2_t(n1778_t),
    .Q(n4697),
    .Q_t(n4697_t)
  );


  nnd2s3
  U3865
  (
    .DIN1(DATA_0_17),
    .DIN1_t(DATA_0_17_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4696),
    .Q_t(n4696_t)
  );


  nnd2s3
  U3866
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1743),
    .DIN2_t(n1743_t),
    .Q(n4695),
    .Q_t(n4695_t)
  );


  nnd4s2
  U3867
  (
    .DIN1(n4702),
    .DIN1_t(n4702_t),
    .DIN2(n4703),
    .DIN2_t(n4703_t),
    .DIN3(n4704),
    .DIN3_t(n4704_t),
    .DIN4(n4705),
    .DIN4_t(n4705_t),
    .Q(WX11014),
    .Q_t(WX11014_t)
  );


  nnd2s3
  U3868
  (
    .DIN1(n2425),
    .DIN1_t(n2425_t),
    .DIN2(n6668),
    .DIN2_t(n6668_t),
    .Q(n4705),
    .Q_t(n4705_t)
  );


  xor2s3
  U3869
  (
    .DIN1(n4706),
    .DIN1_t(n4706_t),
    .DIN2(n4707),
    .DIN2_t(n4707_t),
    .Q(n2425),
    .Q_t(n2425_t)
  );


  xor2s3
  U3870
  (
    .DIN1(n6273),
    .DIN1_t(n6273_t),
    .DIN2(n4708),
    .DIN2_t(n4708_t),
    .Q(n4707),
    .Q_t(n4707_t)
  );


  xor2s3
  U3871
  (
    .DIN1(n6271),
    .DIN1_t(n6271_t),
    .DIN2(n6272),
    .DIN2_t(n6272_t),
    .Q(n4708),
    .Q_t(n4708_t)
  );


  xor2s3
  U3872
  (
    .DIN1(n6274),
    .DIN1_t(n6274_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4706),
    .Q_t(n4706_t)
  );


  nnd2s3
  U3873
  (
    .DIN1(n6595),
    .DIN1_t(n6595_t),
    .DIN2(n1779),
    .DIN2_t(n1779_t),
    .Q(n4704),
    .Q_t(n4704_t)
  );


  nnd2s3
  U3874
  (
    .DIN1(DATA_0_18),
    .DIN1_t(DATA_0_18_t),
    .DIN2(n6637),
    .DIN2_t(n6637_t),
    .Q(n4703),
    .Q_t(n4703_t)
  );


  nnd2s3
  U3875
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n1742),
    .DIN2_t(n1742_t),
    .Q(n4702),
    .Q_t(n4702_t)
  );


  nnd4s2
  U3876
  (
    .DIN1(n4709),
    .DIN1_t(n4709_t),
    .DIN2(n4710),
    .DIN2_t(n4710_t),
    .DIN3(n4711),
    .DIN3_t(n4711_t),
    .DIN4(n4712),
    .DIN4_t(n4712_t),
    .Q(WX11012),
    .Q_t(WX11012_t)
  );


  nnd2s3
  U3877
  (
    .DIN1(n2431),
    .DIN1_t(n2431_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n4712),
    .Q_t(n4712_t)
  );


  xor2s3
  U3878
  (
    .DIN1(n4713),
    .DIN1_t(n4713_t),
    .DIN2(n4714),
    .DIN2_t(n4714_t),
    .Q(n2431),
    .Q_t(n2431_t)
  );


  xor2s3
  U3879
  (
    .DIN1(n6278),
    .DIN1_t(n6278_t),
    .DIN2(n4715),
    .DIN2_t(n4715_t),
    .Q(n4714),
    .Q_t(n4714_t)
  );


  xor2s3
  U3880
  (
    .DIN1(n6276),
    .DIN1_t(n6276_t),
    .DIN2(n6277),
    .DIN2_t(n6277_t),
    .Q(n4715),
    .Q_t(n4715_t)
  );


  xor2s3
  U3881
  (
    .DIN1(n6279),
    .DIN1_t(n6279_t),
    .DIN2(n6695),
    .DIN2_t(n6695_t),
    .Q(n4713),
    .Q_t(n4713_t)
  );


  nnd2s3
  U3882
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1780),
    .DIN2_t(n1780_t),
    .Q(n4711),
    .Q_t(n4711_t)
  );


  nnd2s3
  U3883
  (
    .DIN1(DATA_0_19),
    .DIN1_t(DATA_0_19_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n4710),
    .Q_t(n4710_t)
  );


  nnd2s3
  U3884
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1741),
    .DIN2_t(n1741_t),
    .Q(n4709),
    .Q_t(n4709_t)
  );


  nnd4s2
  U3885
  (
    .DIN1(n4716),
    .DIN1_t(n4716_t),
    .DIN2(n4717),
    .DIN2_t(n4717_t),
    .DIN3(n4718),
    .DIN3_t(n4718_t),
    .DIN4(n4719),
    .DIN4_t(n4719_t),
    .Q(WX11010),
    .Q_t(WX11010_t)
  );


  nnd2s3
  U3886
  (
    .DIN1(n2437),
    .DIN1_t(n2437_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n4719),
    .Q_t(n4719_t)
  );


  xor2s3
  U3887
  (
    .DIN1(n4720),
    .DIN1_t(n4720_t),
    .DIN2(n4721),
    .DIN2_t(n4721_t),
    .Q(n2437),
    .Q_t(n2437_t)
  );


  xor2s3
  U3888
  (
    .DIN1(n6283),
    .DIN1_t(n6283_t),
    .DIN2(n4722),
    .DIN2_t(n4722_t),
    .Q(n4721),
    .Q_t(n4721_t)
  );


  xor2s3
  U3889
  (
    .DIN1(n6281),
    .DIN1_t(n6281_t),
    .DIN2(n6282),
    .DIN2_t(n6282_t),
    .Q(n4722),
    .Q_t(n4722_t)
  );


  xor2s3
  U3890
  (
    .DIN1(n6284),
    .DIN1_t(n6284_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4720),
    .Q_t(n4720_t)
  );


  nnd2s3
  U3891
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1781),
    .DIN2_t(n1781_t),
    .Q(n4718),
    .Q_t(n4718_t)
  );


  nnd2s3
  U3892
  (
    .DIN1(DATA_0_20),
    .DIN1_t(DATA_0_20_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n4717),
    .Q_t(n4717_t)
  );


  nnd2s3
  U3893
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1740),
    .DIN2_t(n1740_t),
    .Q(n4716),
    .Q_t(n4716_t)
  );


  nnd4s2
  U3894
  (
    .DIN1(n4723),
    .DIN1_t(n4723_t),
    .DIN2(n4724),
    .DIN2_t(n4724_t),
    .DIN3(n4725),
    .DIN3_t(n4725_t),
    .DIN4(n4726),
    .DIN4_t(n4726_t),
    .Q(WX11008),
    .Q_t(WX11008_t)
  );


  nnd2s3
  U3895
  (
    .DIN1(n2443),
    .DIN1_t(n2443_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n4726),
    .Q_t(n4726_t)
  );


  xor2s3
  U3896
  (
    .DIN1(n4727),
    .DIN1_t(n4727_t),
    .DIN2(n4728),
    .DIN2_t(n4728_t),
    .Q(n2443),
    .Q_t(n2443_t)
  );


  xor2s3
  U3897
  (
    .DIN1(n6289),
    .DIN1_t(n6289_t),
    .DIN2(n4729),
    .DIN2_t(n4729_t),
    .Q(n4728),
    .Q_t(n4728_t)
  );


  xor2s3
  U3898
  (
    .DIN1(n6287),
    .DIN1_t(n6287_t),
    .DIN2(n6288),
    .DIN2_t(n6288_t),
    .Q(n4729),
    .Q_t(n4729_t)
  );


  xor2s3
  U3899
  (
    .DIN1(n6290),
    .DIN1_t(n6290_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4727),
    .Q_t(n4727_t)
  );


  nnd2s3
  U3900
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1782),
    .DIN2_t(n1782_t),
    .Q(n4725),
    .Q_t(n4725_t)
  );


  nnd2s3
  U3901
  (
    .DIN1(DATA_0_21),
    .DIN1_t(DATA_0_21_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n4724),
    .Q_t(n4724_t)
  );


  nnd2s3
  U3902
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1739),
    .DIN2_t(n1739_t),
    .Q(n4723),
    .Q_t(n4723_t)
  );


  nnd4s2
  U3903
  (
    .DIN1(n4730),
    .DIN1_t(n4730_t),
    .DIN2(n4731),
    .DIN2_t(n4731_t),
    .DIN3(n4732),
    .DIN3_t(n4732_t),
    .DIN4(n4733),
    .DIN4_t(n4733_t),
    .Q(WX11006),
    .Q_t(WX11006_t)
  );


  nnd2s3
  U3904
  (
    .DIN1(n2449),
    .DIN1_t(n2449_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n4733),
    .Q_t(n4733_t)
  );


  xor2s3
  U3905
  (
    .DIN1(n4734),
    .DIN1_t(n4734_t),
    .DIN2(n4735),
    .DIN2_t(n4735_t),
    .Q(n2449),
    .Q_t(n2449_t)
  );


  xor2s3
  U3906
  (
    .DIN1(n6294),
    .DIN1_t(n6294_t),
    .DIN2(n4736),
    .DIN2_t(n4736_t),
    .Q(n4735),
    .Q_t(n4735_t)
  );


  xor2s3
  U3907
  (
    .DIN1(n6292),
    .DIN1_t(n6292_t),
    .DIN2(n6293),
    .DIN2_t(n6293_t),
    .Q(n4736),
    .Q_t(n4736_t)
  );


  xor2s3
  U3908
  (
    .DIN1(n6295),
    .DIN1_t(n6295_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4734),
    .Q_t(n4734_t)
  );


  nnd2s3
  U3909
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1783),
    .DIN2_t(n1783_t),
    .Q(n4732),
    .Q_t(n4732_t)
  );


  nnd2s3
  U3910
  (
    .DIN1(DATA_0_22),
    .DIN1_t(DATA_0_22_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n4731),
    .Q_t(n4731_t)
  );


  nnd2s3
  U3911
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1738),
    .DIN2_t(n1738_t),
    .Q(n4730),
    .Q_t(n4730_t)
  );


  nnd4s2
  U3912
  (
    .DIN1(n4737),
    .DIN1_t(n4737_t),
    .DIN2(n4738),
    .DIN2_t(n4738_t),
    .DIN3(n4739),
    .DIN3_t(n4739_t),
    .DIN4(n4740),
    .DIN4_t(n4740_t),
    .Q(WX11004),
    .Q_t(WX11004_t)
  );


  nnd2s3
  U3913
  (
    .DIN1(n2455),
    .DIN1_t(n2455_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n4740),
    .Q_t(n4740_t)
  );


  xor2s3
  U3914
  (
    .DIN1(n4741),
    .DIN1_t(n4741_t),
    .DIN2(n4742),
    .DIN2_t(n4742_t),
    .Q(n2455),
    .Q_t(n2455_t)
  );


  xor2s3
  U3915
  (
    .DIN1(n6299),
    .DIN1_t(n6299_t),
    .DIN2(n4743),
    .DIN2_t(n4743_t),
    .Q(n4742),
    .Q_t(n4742_t)
  );


  xor2s3
  U3916
  (
    .DIN1(n6297),
    .DIN1_t(n6297_t),
    .DIN2(n6298),
    .DIN2_t(n6298_t),
    .Q(n4743),
    .Q_t(n4743_t)
  );


  xor2s3
  U3917
  (
    .DIN1(n6300),
    .DIN1_t(n6300_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4741),
    .Q_t(n4741_t)
  );


  nnd2s3
  U3918
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1784),
    .DIN2_t(n1784_t),
    .Q(n4739),
    .Q_t(n4739_t)
  );


  nnd2s3
  U3919
  (
    .DIN1(DATA_0_23),
    .DIN1_t(DATA_0_23_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n4738),
    .Q_t(n4738_t)
  );


  nnd2s3
  U3920
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1737),
    .DIN2_t(n1737_t),
    .Q(n4737),
    .Q_t(n4737_t)
  );


  nnd4s2
  U3921
  (
    .DIN1(n4744),
    .DIN1_t(n4744_t),
    .DIN2(n4745),
    .DIN2_t(n4745_t),
    .DIN3(n4746),
    .DIN3_t(n4746_t),
    .DIN4(n4747),
    .DIN4_t(n4747_t),
    .Q(WX11002),
    .Q_t(WX11002_t)
  );


  nnd2s3
  U3922
  (
    .DIN1(n2461),
    .DIN1_t(n2461_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n4747),
    .Q_t(n4747_t)
  );


  xor2s3
  U3923
  (
    .DIN1(n4748),
    .DIN1_t(n4748_t),
    .DIN2(n4749),
    .DIN2_t(n4749_t),
    .Q(n2461),
    .Q_t(n2461_t)
  );


  xor2s3
  U3924
  (
    .DIN1(n6304),
    .DIN1_t(n6304_t),
    .DIN2(n4750),
    .DIN2_t(n4750_t),
    .Q(n4749),
    .Q_t(n4749_t)
  );


  xor2s3
  U3925
  (
    .DIN1(n6302),
    .DIN1_t(n6302_t),
    .DIN2(n6303),
    .DIN2_t(n6303_t),
    .Q(n4750),
    .Q_t(n4750_t)
  );


  xor2s3
  U3926
  (
    .DIN1(n6305),
    .DIN1_t(n6305_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4748),
    .Q_t(n4748_t)
  );


  nnd2s3
  U3927
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1785),
    .DIN2_t(n1785_t),
    .Q(n4746),
    .Q_t(n4746_t)
  );


  nnd2s3
  U3928
  (
    .DIN1(DATA_0_24),
    .DIN1_t(DATA_0_24_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n4745),
    .Q_t(n4745_t)
  );


  nnd2s3
  U3929
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1736),
    .DIN2_t(n1736_t),
    .Q(n4744),
    .Q_t(n4744_t)
  );


  nnd4s2
  U3930
  (
    .DIN1(n4751),
    .DIN1_t(n4751_t),
    .DIN2(n4752),
    .DIN2_t(n4752_t),
    .DIN3(n4753),
    .DIN3_t(n4753_t),
    .DIN4(n4754),
    .DIN4_t(n4754_t),
    .Q(WX11000),
    .Q_t(WX11000_t)
  );


  nnd2s3
  U3931
  (
    .DIN1(n2467),
    .DIN1_t(n2467_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n4754),
    .Q_t(n4754_t)
  );


  xor2s3
  U3932
  (
    .DIN1(n4755),
    .DIN1_t(n4755_t),
    .DIN2(n4756),
    .DIN2_t(n4756_t),
    .Q(n2467),
    .Q_t(n2467_t)
  );


  xor2s3
  U3933
  (
    .DIN1(n6309),
    .DIN1_t(n6309_t),
    .DIN2(n4757),
    .DIN2_t(n4757_t),
    .Q(n4756),
    .Q_t(n4756_t)
  );


  xor2s3
  U3934
  (
    .DIN1(n6307),
    .DIN1_t(n6307_t),
    .DIN2(n6308),
    .DIN2_t(n6308_t),
    .Q(n4757),
    .Q_t(n4757_t)
  );


  xor2s3
  U3935
  (
    .DIN1(n6310),
    .DIN1_t(n6310_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4755),
    .Q_t(n4755_t)
  );


  nnd2s3
  U3936
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1786),
    .DIN2_t(n1786_t),
    .Q(n4753),
    .Q_t(n4753_t)
  );


  nnd2s3
  U3937
  (
    .DIN1(DATA_0_25),
    .DIN1_t(DATA_0_25_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n4752),
    .Q_t(n4752_t)
  );


  nnd2s3
  U3938
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1735),
    .DIN2_t(n1735_t),
    .Q(n4751),
    .Q_t(n4751_t)
  );


  nnd4s2
  U3939
  (
    .DIN1(n4758),
    .DIN1_t(n4758_t),
    .DIN2(n4759),
    .DIN2_t(n4759_t),
    .DIN3(n4760),
    .DIN3_t(n4760_t),
    .DIN4(n4761),
    .DIN4_t(n4761_t),
    .Q(WX10998),
    .Q_t(WX10998_t)
  );


  nnd2s3
  U3940
  (
    .DIN1(n2473),
    .DIN1_t(n2473_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n4761),
    .Q_t(n4761_t)
  );


  xor2s3
  U3941
  (
    .DIN1(n4762),
    .DIN1_t(n4762_t),
    .DIN2(n4763),
    .DIN2_t(n4763_t),
    .Q(n2473),
    .Q_t(n2473_t)
  );


  xor2s3
  U3942
  (
    .DIN1(n6314),
    .DIN1_t(n6314_t),
    .DIN2(n4764),
    .DIN2_t(n4764_t),
    .Q(n4763),
    .Q_t(n4763_t)
  );


  xor2s3
  U3943
  (
    .DIN1(n6312),
    .DIN1_t(n6312_t),
    .DIN2(n6313),
    .DIN2_t(n6313_t),
    .Q(n4764),
    .Q_t(n4764_t)
  );


  xor2s3
  U3944
  (
    .DIN1(n6315),
    .DIN1_t(n6315_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4762),
    .Q_t(n4762_t)
  );


  nnd2s3
  U3945
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1787),
    .DIN2_t(n1787_t),
    .Q(n4760),
    .Q_t(n4760_t)
  );


  nnd2s3
  U3946
  (
    .DIN1(DATA_0_26),
    .DIN1_t(DATA_0_26_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n4759),
    .Q_t(n4759_t)
  );


  nnd2s3
  U3947
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1734),
    .DIN2_t(n1734_t),
    .Q(n4758),
    .Q_t(n4758_t)
  );


  nnd4s2
  U3948
  (
    .DIN1(n4765),
    .DIN1_t(n4765_t),
    .DIN2(n4766),
    .DIN2_t(n4766_t),
    .DIN3(n4767),
    .DIN3_t(n4767_t),
    .DIN4(n4768),
    .DIN4_t(n4768_t),
    .Q(WX10996),
    .Q_t(WX10996_t)
  );


  nnd2s3
  U3949
  (
    .DIN1(n2479),
    .DIN1_t(n2479_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n4768),
    .Q_t(n4768_t)
  );


  xor2s3
  U3950
  (
    .DIN1(n4769),
    .DIN1_t(n4769_t),
    .DIN2(n4770),
    .DIN2_t(n4770_t),
    .Q(n2479),
    .Q_t(n2479_t)
  );


  xor2s3
  U3951
  (
    .DIN1(n6319),
    .DIN1_t(n6319_t),
    .DIN2(n4771),
    .DIN2_t(n4771_t),
    .Q(n4770),
    .Q_t(n4770_t)
  );


  xor2s3
  U3952
  (
    .DIN1(n6317),
    .DIN1_t(n6317_t),
    .DIN2(n6318),
    .DIN2_t(n6318_t),
    .Q(n4771),
    .Q_t(n4771_t)
  );


  xor2s3
  U3953
  (
    .DIN1(n6320),
    .DIN1_t(n6320_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4769),
    .Q_t(n4769_t)
  );


  nnd2s3
  U3954
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1788),
    .DIN2_t(n1788_t),
    .Q(n4767),
    .Q_t(n4767_t)
  );


  nnd2s3
  U3955
  (
    .DIN1(DATA_0_27),
    .DIN1_t(DATA_0_27_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n4766),
    .Q_t(n4766_t)
  );


  nnd2s3
  U3956
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1733),
    .DIN2_t(n1733_t),
    .Q(n4765),
    .Q_t(n4765_t)
  );


  nnd4s2
  U3957
  (
    .DIN1(n4772),
    .DIN1_t(n4772_t),
    .DIN2(n4773),
    .DIN2_t(n4773_t),
    .DIN3(n4774),
    .DIN3_t(n4774_t),
    .DIN4(n4775),
    .DIN4_t(n4775_t),
    .Q(WX10994),
    .Q_t(WX10994_t)
  );


  nnd2s3
  U3958
  (
    .DIN1(n2485),
    .DIN1_t(n2485_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n4775),
    .Q_t(n4775_t)
  );


  xor2s3
  U3959
  (
    .DIN1(n4776),
    .DIN1_t(n4776_t),
    .DIN2(n4777),
    .DIN2_t(n4777_t),
    .Q(n2485),
    .Q_t(n2485_t)
  );


  xor2s3
  U3960
  (
    .DIN1(n6324),
    .DIN1_t(n6324_t),
    .DIN2(n4778),
    .DIN2_t(n4778_t),
    .Q(n4777),
    .Q_t(n4777_t)
  );


  xor2s3
  U3961
  (
    .DIN1(n6322),
    .DIN1_t(n6322_t),
    .DIN2(n6323),
    .DIN2_t(n6323_t),
    .Q(n4778),
    .Q_t(n4778_t)
  );


  xor2s3
  U3962
  (
    .DIN1(n6325),
    .DIN1_t(n6325_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4776),
    .Q_t(n4776_t)
  );


  nnd2s3
  U3963
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1789),
    .DIN2_t(n1789_t),
    .Q(n4774),
    .Q_t(n4774_t)
  );


  nnd2s3
  U3964
  (
    .DIN1(DATA_0_28),
    .DIN1_t(DATA_0_28_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n4773),
    .Q_t(n4773_t)
  );


  nnd2s3
  U3965
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1732),
    .DIN2_t(n1732_t),
    .Q(n4772),
    .Q_t(n4772_t)
  );


  nnd4s2
  U3966
  (
    .DIN1(n4779),
    .DIN1_t(n4779_t),
    .DIN2(n4780),
    .DIN2_t(n4780_t),
    .DIN3(n4781),
    .DIN3_t(n4781_t),
    .DIN4(n4782),
    .DIN4_t(n4782_t),
    .Q(WX10992),
    .Q_t(WX10992_t)
  );


  nnd2s3
  U3967
  (
    .DIN1(n2491),
    .DIN1_t(n2491_t),
    .DIN2(n6667),
    .DIN2_t(n6667_t),
    .Q(n4782),
    .Q_t(n4782_t)
  );


  xor2s3
  U3968
  (
    .DIN1(n4783),
    .DIN1_t(n4783_t),
    .DIN2(n4784),
    .DIN2_t(n4784_t),
    .Q(n2491),
    .Q_t(n2491_t)
  );


  xor2s3
  U3969
  (
    .DIN1(n6329),
    .DIN1_t(n6329_t),
    .DIN2(n4785),
    .DIN2_t(n4785_t),
    .Q(n4784),
    .Q_t(n4784_t)
  );


  xor2s3
  U3970
  (
    .DIN1(n6327),
    .DIN1_t(n6327_t),
    .DIN2(n6328),
    .DIN2_t(n6328_t),
    .Q(n4785),
    .Q_t(n4785_t)
  );


  xor2s3
  U3971
  (
    .DIN1(n6330),
    .DIN1_t(n6330_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4783),
    .Q_t(n4783_t)
  );


  nnd2s3
  U3972
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1790),
    .DIN2_t(n1790_t),
    .Q(n4781),
    .Q_t(n4781_t)
  );


  nnd2s3
  U3973
  (
    .DIN1(DATA_0_29),
    .DIN1_t(DATA_0_29_t),
    .DIN2(n6636),
    .DIN2_t(n6636_t),
    .Q(n4780),
    .Q_t(n4780_t)
  );


  nnd2s3
  U3974
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1731),
    .DIN2_t(n1731_t),
    .Q(n4779),
    .Q_t(n4779_t)
  );


  nnd4s2
  U3975
  (
    .DIN1(n4786),
    .DIN1_t(n4786_t),
    .DIN2(n4787),
    .DIN2_t(n4787_t),
    .DIN3(n4788),
    .DIN3_t(n4788_t),
    .DIN4(n4789),
    .DIN4_t(n4789_t),
    .Q(WX10990),
    .Q_t(WX10990_t)
  );


  nnd2s3
  U3976
  (
    .DIN1(n2497),
    .DIN1_t(n2497_t),
    .DIN2(n6672),
    .DIN2_t(n6672_t),
    .Q(n4789),
    .Q_t(n4789_t)
  );


  xor2s3
  U3977
  (
    .DIN1(n4790),
    .DIN1_t(n4790_t),
    .DIN2(n4791),
    .DIN2_t(n4791_t),
    .Q(n2497),
    .Q_t(n2497_t)
  );


  xor2s3
  U3978
  (
    .DIN1(n6334),
    .DIN1_t(n6334_t),
    .DIN2(n4792),
    .DIN2_t(n4792_t),
    .Q(n4791),
    .Q_t(n4791_t)
  );


  xor2s3
  U3979
  (
    .DIN1(n6332),
    .DIN1_t(n6332_t),
    .DIN2(n6333),
    .DIN2_t(n6333_t),
    .Q(n4792),
    .Q_t(n4792_t)
  );


  xor2s3
  U3980
  (
    .DIN1(n6335),
    .DIN1_t(n6335_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4790),
    .Q_t(n4790_t)
  );


  nnd2s3
  U3981
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1791),
    .DIN2_t(n1791_t),
    .Q(n4788),
    .Q_t(n4788_t)
  );


  nnd2s3
  U3982
  (
    .DIN1(DATA_0_30),
    .DIN1_t(DATA_0_30_t),
    .DIN2(n6641),
    .DIN2_t(n6641_t),
    .Q(n4787),
    .Q_t(n4787_t)
  );


  nnd2s3
  U3983
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1730),
    .DIN2_t(n1730_t),
    .Q(n4786),
    .Q_t(n4786_t)
  );


  nnd4s2
  U3984
  (
    .DIN1(n4793),
    .DIN1_t(n4793_t),
    .DIN2(n4794),
    .DIN2_t(n4794_t),
    .DIN3(n4795),
    .DIN3_t(n4795_t),
    .DIN4(n4796),
    .DIN4_t(n4796_t),
    .Q(WX10988),
    .Q_t(WX10988_t)
  );


  nnd2s3
  U3985
  (
    .DIN1(n6594),
    .DIN1_t(n6594_t),
    .DIN2(n1792),
    .DIN2_t(n1792_t),
    .Q(n4796),
    .Q_t(n4796_t)
  );


  and3s3
  U3986
  (
    .DIN1(TM1),
    .DIN1_t(TM1_t),
    .DIN2(RESET),
    .DIN2_t(RESET_t),
    .DIN3(n6703),
    .DIN3_t(n6703_t),
    .Q(n2316),
    .Q_t(n2316_t)
  );


  nnd2s3
  U3987
  (
    .DIN1(DATA_0_31),
    .DIN1_t(DATA_0_31_t),
    .DIN2(n6625),
    .DIN2_t(n6625_t),
    .Q(n4795),
    .Q_t(n4795_t)
  );


  and3s3
  U3988
  (
    .DIN1(n6711),
    .DIN1_t(n6711_t),
    .DIN2(n6698),
    .DIN2_t(n6698_t),
    .DIN3(RESET),
    .DIN3_t(RESET_t),
    .Q(n2314),
    .Q_t(n2314_t)
  );


  nnd2s3
  U3989
  (
    .DIN1(n6563),
    .DIN1_t(n6563_t),
    .DIN2(n1729),
    .DIN2_t(n1729_t),
    .Q(n4794),
    .Q_t(n4794_t)
  );


  and3s3
  U3990
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6698),
    .DIN2_t(n6698_t),
    .DIN3(n6703),
    .DIN3_t(n6703_t),
    .Q(n2317),
    .Q_t(n2317_t)
  );


  nnd2s3
  U3991
  (
    .DIN1(n2503),
    .DIN1_t(n2503_t),
    .DIN2(n6661),
    .DIN2_t(n6661_t),
    .Q(n4793),
    .Q_t(n4793_t)
  );


  and3s3
  U3992
  (
    .DIN1(RESET),
    .DIN1_t(RESET_t),
    .DIN2(n6711),
    .DIN2_t(n6711_t),
    .DIN3(TM1),
    .DIN3_t(TM1_t),
    .Q(n2312),
    .Q_t(n2312_t)
  );


  xor2s3
  U3993
  (
    .DIN1(n4797),
    .DIN1_t(n4797_t),
    .DIN2(n4798),
    .DIN2_t(n4798_t),
    .Q(n2503),
    .Q_t(n2503_t)
  );


  xor2s3
  U3994
  (
    .DIN1(n6340),
    .DIN1_t(n6340_t),
    .DIN2(n4799),
    .DIN2_t(n4799_t),
    .Q(n4798),
    .Q_t(n4798_t)
  );


  xor2s3
  U3995
  (
    .DIN1(n6338),
    .DIN1_t(n6338_t),
    .DIN2(n6339),
    .DIN2_t(n6339_t),
    .Q(n4799),
    .Q_t(n4799_t)
  );


  xor2s3
  U3996
  (
    .DIN1(n6341),
    .DIN1_t(n6341_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4797),
    .Q_t(n4797_t)
  );


  nor2s3
  U3997
  (
    .DIN1(n6789),
    .DIN1_t(n6789_t),
    .DIN2(n1792),
    .DIN2_t(n1792_t),
    .Q(WX10890),
    .Q_t(WX10890_t)
  );


  nor2s3
  U3998
  (
    .DIN1(n6344),
    .DIN1_t(n6344_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX10888),
    .Q_t(WX10888_t)
  );


  nor2s3
  U3999
  (
    .DIN1(n6345),
    .DIN1_t(n6345_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX10886),
    .Q_t(WX10886_t)
  );


  nor2s3
  U4000
  (
    .DIN1(n6346),
    .DIN1_t(n6346_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX10884),
    .Q_t(WX10884_t)
  );


  nor2s3
  U4001
  (
    .DIN1(n6347),
    .DIN1_t(n6347_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX10882),
    .Q_t(WX10882_t)
  );


  nor2s3
  U4002
  (
    .DIN1(n6348),
    .DIN1_t(n6348_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX10880),
    .Q_t(WX10880_t)
  );


  nor2s3
  U4003
  (
    .DIN1(n6349),
    .DIN1_t(n6349_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX10878),
    .Q_t(WX10878_t)
  );


  nor2s3
  U4004
  (
    .DIN1(n6350),
    .DIN1_t(n6350_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX10876),
    .Q_t(WX10876_t)
  );


  nor2s3
  U4005
  (
    .DIN1(n6351),
    .DIN1_t(n6351_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX10874),
    .Q_t(WX10874_t)
  );


  nor2s3
  U4006
  (
    .DIN1(n6352),
    .DIN1_t(n6352_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX10872),
    .Q_t(WX10872_t)
  );


  nor2s3
  U4007
  (
    .DIN1(n6353),
    .DIN1_t(n6353_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX10870),
    .Q_t(WX10870_t)
  );


  nor2s3
  U4008
  (
    .DIN1(n6355),
    .DIN1_t(n6355_t),
    .DIN2(n6768),
    .DIN2_t(n6768_t),
    .Q(WX10868),
    .Q_t(WX10868_t)
  );


  nor2s3
  U4009
  (
    .DIN1(n6356),
    .DIN1_t(n6356_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10866),
    .Q_t(WX10866_t)
  );


  nor2s3
  U4010
  (
    .DIN1(n6357),
    .DIN1_t(n6357_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10864),
    .Q_t(WX10864_t)
  );


  nor2s3
  U4011
  (
    .DIN1(n6358),
    .DIN1_t(n6358_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10862),
    .Q_t(WX10862_t)
  );


  nor2s3
  U4012
  (
    .DIN1(n6359),
    .DIN1_t(n6359_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10860),
    .Q_t(WX10860_t)
  );


  nor2s3
  U4013
  (
    .DIN1(n6360),
    .DIN1_t(n6360_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10858),
    .Q_t(WX10858_t)
  );


  nor2s3
  U4014
  (
    .DIN1(n6361),
    .DIN1_t(n6361_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10856),
    .Q_t(WX10856_t)
  );


  nor2s3
  U4015
  (
    .DIN1(n6362),
    .DIN1_t(n6362_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10854),
    .Q_t(WX10854_t)
  );


  nor2s3
  U4016
  (
    .DIN1(n6363),
    .DIN1_t(n6363_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10852),
    .Q_t(WX10852_t)
  );


  nor2s3
  U4017
  (
    .DIN1(n6364),
    .DIN1_t(n6364_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10850),
    .Q_t(WX10850_t)
  );


  nor2s3
  U4018
  (
    .DIN1(n6365),
    .DIN1_t(n6365_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10848),
    .Q_t(WX10848_t)
  );


  nor2s3
  U4019
  (
    .DIN1(n6366),
    .DIN1_t(n6366_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10846),
    .Q_t(WX10846_t)
  );


  nor2s3
  U4020
  (
    .DIN1(n6367),
    .DIN1_t(n6367_t),
    .DIN2(n6767),
    .DIN2_t(n6767_t),
    .Q(WX10844),
    .Q_t(WX10844_t)
  );


  nor2s3
  U4021
  (
    .DIN1(n6368),
    .DIN1_t(n6368_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX10842),
    .Q_t(WX10842_t)
  );


  nor2s3
  U4022
  (
    .DIN1(n6369),
    .DIN1_t(n6369_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX10840),
    .Q_t(WX10840_t)
  );


  nor2s3
  U4023
  (
    .DIN1(n6370),
    .DIN1_t(n6370_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX10838),
    .Q_t(WX10838_t)
  );


  nor2s3
  U4024
  (
    .DIN1(n6371),
    .DIN1_t(n6371_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX10836),
    .Q_t(WX10836_t)
  );


  nor2s3
  U4025
  (
    .DIN1(n6372),
    .DIN1_t(n6372_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX10834),
    .Q_t(WX10834_t)
  );


  nor2s3
  U4026
  (
    .DIN1(n6373),
    .DIN1_t(n6373_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX10832),
    .Q_t(WX10832_t)
  );


  nor2s3
  U4027
  (
    .DIN1(n6374),
    .DIN1_t(n6374_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX10830),
    .Q_t(WX10830_t)
  );


  nor2s3
  U4028
  (
    .DIN1(n6375),
    .DIN1_t(n6375_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX10828),
    .Q_t(WX10828_t)
  );


  nor2s3
  U4029
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n4800),
    .DIN2_t(n4800_t),
    .Q(WX10377),
    .Q_t(WX10377_t)
  );


  xor2s3
  U4030
  (
    .DIN1(n6383),
    .DIN1_t(n6383_t),
    .DIN2(n6384),
    .DIN2_t(n6384_t),
    .Q(n4800),
    .Q_t(n4800_t)
  );


  nor2s3
  U4031
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n4801),
    .DIN2_t(n4801_t),
    .Q(WX10375),
    .Q_t(WX10375_t)
  );


  xor2s3
  U4032
  (
    .DIN1(n6385),
    .DIN1_t(n6385_t),
    .DIN2(n6386),
    .DIN2_t(n6386_t),
    .Q(n4801),
    .Q_t(n4801_t)
  );


  nor2s3
  U4033
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n4802),
    .DIN2_t(n4802_t),
    .Q(WX10373),
    .Q_t(WX10373_t)
  );


  xor2s3
  U4034
  (
    .DIN1(n6387),
    .DIN1_t(n6387_t),
    .DIN2(n6388),
    .DIN2_t(n6388_t),
    .Q(n4802),
    .Q_t(n4802_t)
  );


  nor2s3
  U4035
  (
    .DIN1(n6795),
    .DIN1_t(n6795_t),
    .DIN2(n4803),
    .DIN2_t(n4803_t),
    .Q(WX10371),
    .Q_t(WX10371_t)
  );


  xor2s3
  U4036
  (
    .DIN1(n6389),
    .DIN1_t(n6389_t),
    .DIN2(n6390),
    .DIN2_t(n6390_t),
    .Q(n4803),
    .Q_t(n4803_t)
  );


  nor2s3
  U4037
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n4804),
    .DIN2_t(n4804_t),
    .Q(WX10369),
    .Q_t(WX10369_t)
  );


  xor2s3
  U4038
  (
    .DIN1(n6391),
    .DIN1_t(n6391_t),
    .DIN2(n6392),
    .DIN2_t(n6392_t),
    .Q(n4804),
    .Q_t(n4804_t)
  );


  nor2s3
  U4039
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n4805),
    .DIN2_t(n4805_t),
    .Q(WX10367),
    .Q_t(WX10367_t)
  );


  xor2s3
  U4040
  (
    .DIN1(n6393),
    .DIN1_t(n6393_t),
    .DIN2(n6394),
    .DIN2_t(n6394_t),
    .Q(n4805),
    .Q_t(n4805_t)
  );


  nor2s3
  U4041
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n4806),
    .DIN2_t(n4806_t),
    .Q(WX10365),
    .Q_t(WX10365_t)
  );


  xor2s3
  U4042
  (
    .DIN1(n6395),
    .DIN1_t(n6395_t),
    .DIN2(n6396),
    .DIN2_t(n6396_t),
    .Q(n4806),
    .Q_t(n4806_t)
  );


  nor2s3
  U4043
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n4807),
    .DIN2_t(n4807_t),
    .Q(WX10363),
    .Q_t(WX10363_t)
  );


  xor2s3
  U4044
  (
    .DIN1(n6397),
    .DIN1_t(n6397_t),
    .DIN2(n6398),
    .DIN2_t(n6398_t),
    .Q(n4807),
    .Q_t(n4807_t)
  );


  nor2s3
  U4045
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n4808),
    .DIN2_t(n4808_t),
    .Q(WX10361),
    .Q_t(WX10361_t)
  );


  xor2s3
  U4046
  (
    .DIN1(n6399),
    .DIN1_t(n6399_t),
    .DIN2(n6400),
    .DIN2_t(n6400_t),
    .Q(n4808),
    .Q_t(n4808_t)
  );


  nor2s3
  U4047
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n4809),
    .DIN2_t(n4809_t),
    .Q(WX10359),
    .Q_t(WX10359_t)
  );


  xor2s3
  U4048
  (
    .DIN1(n6401),
    .DIN1_t(n6401_t),
    .DIN2(n6402),
    .DIN2_t(n6402_t),
    .Q(n4809),
    .Q_t(n4809_t)
  );


  nor2s3
  U4049
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n4810),
    .DIN2_t(n4810_t),
    .Q(WX10357),
    .Q_t(WX10357_t)
  );


  xor2s3
  U4050
  (
    .DIN1(n6403),
    .DIN1_t(n6403_t),
    .DIN2(n6404),
    .DIN2_t(n6404_t),
    .Q(n4810),
    .Q_t(n4810_t)
  );


  nor2s3
  U4051
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n4811),
    .DIN2_t(n4811_t),
    .Q(WX10355),
    .Q_t(WX10355_t)
  );


  xor2s3
  U4052
  (
    .DIN1(n6405),
    .DIN1_t(n6405_t),
    .DIN2(n6406),
    .DIN2_t(n6406_t),
    .Q(n4811),
    .Q_t(n4811_t)
  );


  nor2s3
  U4053
  (
    .DIN1(n6794),
    .DIN1_t(n6794_t),
    .DIN2(n4812),
    .DIN2_t(n4812_t),
    .Q(WX10353),
    .Q_t(WX10353_t)
  );


  xor2s3
  U4054
  (
    .DIN1(n6407),
    .DIN1_t(n6407_t),
    .DIN2(n6408),
    .DIN2_t(n6408_t),
    .Q(n4812),
    .Q_t(n4812_t)
  );


  nor2s3
  U4055
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n4813),
    .DIN2_t(n4813_t),
    .Q(WX10351),
    .Q_t(WX10351_t)
  );


  xor2s3
  U4056
  (
    .DIN1(n6409),
    .DIN1_t(n6409_t),
    .DIN2(n6410),
    .DIN2_t(n6410_t),
    .Q(n4813),
    .Q_t(n4813_t)
  );


  nor2s3
  U4057
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n4814),
    .DIN2_t(n4814_t),
    .Q(WX10349),
    .Q_t(WX10349_t)
  );


  xor2s3
  U4058
  (
    .DIN1(n6411),
    .DIN1_t(n6411_t),
    .DIN2(n6412),
    .DIN2_t(n6412_t),
    .Q(n4814),
    .Q_t(n4814_t)
  );


  nor2s3
  U4059
  (
    .DIN1(n4815),
    .DIN1_t(n4815_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX10347),
    .Q_t(WX10347_t)
  );


  xor2s3
  U4060
  (
    .DIN1(n1793),
    .DIN1_t(n1793_t),
    .DIN2(n4816),
    .DIN2_t(n4816_t),
    .Q(n4815),
    .Q_t(n4815_t)
  );


  xor2s3
  U4061
  (
    .DIN1(n6413),
    .DIN1_t(n6413_t),
    .DIN2(n6414),
    .DIN2_t(n6414_t),
    .Q(n4816),
    .Q_t(n4816_t)
  );


  nor2s3
  U4062
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n4817),
    .DIN2_t(n4817_t),
    .Q(WX10345),
    .Q_t(WX10345_t)
  );


  xor2s3
  U4063
  (
    .DIN1(n6415),
    .DIN1_t(n6415_t),
    .DIN2(n3220),
    .DIN2_t(n3220_t),
    .Q(n4817),
    .Q_t(n4817_t)
  );


  nor2s3
  U4064
  (
    .DIN1(n6793),
    .DIN1_t(n6793_t),
    .DIN2(n4818),
    .DIN2_t(n4818_t),
    .Q(WX10343),
    .Q_t(WX10343_t)
  );


  xor2s3
  U4065
  (
    .DIN1(n6416),
    .DIN1_t(n6416_t),
    .DIN2(n3219),
    .DIN2_t(n3219_t),
    .Q(n4818),
    .Q_t(n4818_t)
  );


  nor2s3
  U4066
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n4819),
    .DIN2_t(n4819_t),
    .Q(WX10341),
    .Q_t(WX10341_t)
  );


  xor2s3
  U4067
  (
    .DIN1(n6417),
    .DIN1_t(n6417_t),
    .DIN2(n3218),
    .DIN2_t(n3218_t),
    .Q(n4819),
    .Q_t(n4819_t)
  );


  nor2s3
  U4068
  (
    .DIN1(n6792),
    .DIN1_t(n6792_t),
    .DIN2(n4820),
    .DIN2_t(n4820_t),
    .Q(WX10339),
    .Q_t(WX10339_t)
  );


  xor2s3
  U4069
  (
    .DIN1(n6418),
    .DIN1_t(n6418_t),
    .DIN2(n3217),
    .DIN2_t(n3217_t),
    .Q(n4820),
    .Q_t(n4820_t)
  );


  nor2s3
  U4070
  (
    .DIN1(n4821),
    .DIN1_t(n4821_t),
    .DIN2(n6766),
    .DIN2_t(n6766_t),
    .Q(WX10337),
    .Q_t(WX10337_t)
  );


  xnr2s3
  U4071
  (
    .DIN1(n3216),
    .DIN1_t(n3216_t),
    .DIN2(n4822),
    .DIN2_t(n4822_t),
    .Q(n4821),
    .Q_t(n4821_t)
  );


  xor2s3
  U4072
  (
    .DIN1(n6419),
    .DIN1_t(n6419_t),
    .DIN2(n6430),
    .DIN2_t(n6430_t),
    .Q(n4822),
    .Q_t(n4822_t)
  );


  nor2s3
  U4073
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n4823),
    .DIN2_t(n4823_t),
    .Q(WX10335),
    .Q_t(WX10335_t)
  );


  xor2s3
  U4074
  (
    .DIN1(n6420),
    .DIN1_t(n6420_t),
    .DIN2(n3215),
    .DIN2_t(n3215_t),
    .Q(n4823),
    .Q_t(n4823_t)
  );


  nor2s3
  U4075
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n4824),
    .DIN2_t(n4824_t),
    .Q(WX10333),
    .Q_t(WX10333_t)
  );


  xor2s3
  U4076
  (
    .DIN1(n6421),
    .DIN1_t(n6421_t),
    .DIN2(n3214),
    .DIN2_t(n3214_t),
    .Q(n4824),
    .Q_t(n4824_t)
  );


  nor2s3
  U4077
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n4825),
    .DIN2_t(n4825_t),
    .Q(WX10331),
    .Q_t(WX10331_t)
  );


  xor2s3
  U4078
  (
    .DIN1(n6422),
    .DIN1_t(n6422_t),
    .DIN2(n3213),
    .DIN2_t(n3213_t),
    .Q(n4825),
    .Q_t(n4825_t)
  );


  nor2s3
  U4079
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n4826),
    .DIN2_t(n4826_t),
    .Q(WX10329),
    .Q_t(WX10329_t)
  );


  xor2s3
  U4080
  (
    .DIN1(n6423),
    .DIN1_t(n6423_t),
    .DIN2(n3212),
    .DIN2_t(n3212_t),
    .Q(n4826),
    .Q_t(n4826_t)
  );


  nor2s3
  U4081
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n4827),
    .DIN2_t(n4827_t),
    .Q(WX10327),
    .Q_t(WX10327_t)
  );


  xor2s3
  U4082
  (
    .DIN1(n6424),
    .DIN1_t(n6424_t),
    .DIN2(n3211),
    .DIN2_t(n3211_t),
    .Q(n4827),
    .Q_t(n4827_t)
  );


  nor2s3
  U4083
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n4828),
    .DIN2_t(n4828_t),
    .Q(WX10325),
    .Q_t(WX10325_t)
  );


  xor2s3
  U4084
  (
    .DIN1(n6425),
    .DIN1_t(n6425_t),
    .DIN2(n3210),
    .DIN2_t(n3210_t),
    .Q(n4828),
    .Q_t(n4828_t)
  );


  nor2s3
  U4085
  (
    .DIN1(n4829),
    .DIN1_t(n4829_t),
    .DIN2(n6771),
    .DIN2_t(n6771_t),
    .Q(WX10323),
    .Q_t(WX10323_t)
  );


  xnr2s3
  U4086
  (
    .DIN1(n3209),
    .DIN1_t(n3209_t),
    .DIN2(n4830),
    .DIN2_t(n4830_t),
    .Q(n4829),
    .Q_t(n4829_t)
  );


  xor2s3
  U4087
  (
    .DIN1(n6426),
    .DIN1_t(n6426_t),
    .DIN2(n6430),
    .DIN2_t(n6430_t),
    .Q(n4830),
    .Q_t(n4830_t)
  );


  nor2s3
  U4088
  (
    .DIN1(n6791),
    .DIN1_t(n6791_t),
    .DIN2(n4831),
    .DIN2_t(n4831_t),
    .Q(WX10321),
    .Q_t(WX10321_t)
  );


  xor2s3
  U4089
  (
    .DIN1(n6427),
    .DIN1_t(n6427_t),
    .DIN2(n3208),
    .DIN2_t(n3208_t),
    .Q(n4831),
    .Q_t(n4831_t)
  );


  nor2s3
  U4090
  (
    .DIN1(n6790),
    .DIN1_t(n6790_t),
    .DIN2(n4832),
    .DIN2_t(n4832_t),
    .Q(WX10319),
    .Q_t(WX10319_t)
  );


  xor2s3
  U4091
  (
    .DIN1(n6428),
    .DIN1_t(n6428_t),
    .DIN2(n3207),
    .DIN2_t(n3207_t),
    .Q(n4832),
    .Q_t(n4832_t)
  );


  nor2s3
  U4092
  (
    .DIN1(n6788),
    .DIN1_t(n6788_t),
    .DIN2(n4833),
    .DIN2_t(n4833_t),
    .Q(WX10317),
    .Q_t(WX10317_t)
  );


  xor2s3
  U4093
  (
    .DIN1(n6429),
    .DIN1_t(n6429_t),
    .DIN2(n3206),
    .DIN2_t(n3206_t),
    .Q(n4833),
    .Q_t(n4833_t)
  );


  nor2s3
  U4094
  (
    .DIN1(n6788),
    .DIN1_t(n6788_t),
    .DIN2(n4834),
    .DIN2_t(n4834_t),
    .Q(WX10315),
    .Q_t(WX10315_t)
  );


  xor2s3
  U4095
  (
    .DIN1(n6430),
    .DIN1_t(n6430_t),
    .DIN2(n3205),
    .DIN2_t(n3205_t),
    .Q(n4834),
    .Q_t(n4834_t)
  );


  xnr2s3
  U4096
  (
    .DIN1(n4835),
    .DIN1_t(n4835_t),
    .DIN2(n3113),
    .DIN2_t(n3113_t),
    .Q(DATA_9_9),
    .Q_t(DATA_9_9_t)
  );


  xnr2s3
  U4097
  (
    .DIN1(n4836),
    .DIN1_t(n4836_t),
    .DIN2(n4837),
    .DIN2_t(n4837_t),
    .Q(n3113),
    .Q_t(n3113_t)
  );


  xor2s3
  U4098
  (
    .DIN1(n6506),
    .DIN1_t(n6506_t),
    .DIN2(n4838),
    .DIN2_t(n4838_t),
    .Q(n4837),
    .Q_t(n4837_t)
  );


  xor2s3
  U4099
  (
    .DIN1(n6504),
    .DIN1_t(n6504_t),
    .DIN2(n6505),
    .DIN2_t(n6505_t),
    .Q(n4838),
    .Q_t(n4838_t)
  );


  xor2s3
  U4100
  (
    .DIN1(n6507),
    .DIN1_t(n6507_t),
    .DIN2(n6710),
    .DIN2_t(n6710_t),
    .Q(n4836),
    .Q_t(n4836_t)
  );


  nnd2s3
  U4101
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2282),
    .DIN2_t(n2282_t),
    .Q(n4835),
    .Q_t(n4835_t)
  );


  xnr2s3
  U4102
  (
    .DIN1(n4839),
    .DIN1_t(n4839_t),
    .DIN2(n3107),
    .DIN2_t(n3107_t),
    .Q(DATA_9_8),
    .Q_t(DATA_9_8_t)
  );


  xnr2s3
  U4103
  (
    .DIN1(n4840),
    .DIN1_t(n4840_t),
    .DIN2(n4841),
    .DIN2_t(n4841_t),
    .Q(n3107),
    .Q_t(n3107_t)
  );


  xor2s3
  U4104
  (
    .DIN1(n6455),
    .DIN1_t(n6455_t),
    .DIN2(n4842),
    .DIN2_t(n4842_t),
    .Q(n4841),
    .Q_t(n4841_t)
  );


  xor2s3
  U4105
  (
    .DIN1(n6453),
    .DIN1_t(n6453_t),
    .DIN2(n6454),
    .DIN2_t(n6454_t),
    .Q(n4842),
    .Q_t(n4842_t)
  );


  xor2s3
  U4106
  (
    .DIN1(n6556),
    .DIN1_t(n6556_t),
    .DIN2(n6710),
    .DIN2_t(n6710_t),
    .Q(n4840),
    .Q_t(n4840_t)
  );


  nnd2s3
  U4107
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2281),
    .DIN2_t(n2281_t),
    .Q(n4839),
    .Q_t(n4839_t)
  );


  xnr2s3
  U4108
  (
    .DIN1(n4843),
    .DIN1_t(n4843_t),
    .DIN2(n3101),
    .DIN2_t(n3101_t),
    .Q(DATA_9_7),
    .Q_t(DATA_9_7_t)
  );


  xnr2s3
  U4109
  (
    .DIN1(n4844),
    .DIN1_t(n4844_t),
    .DIN2(n4845),
    .DIN2_t(n4845_t),
    .Q(n3101),
    .Q_t(n3101_t)
  );


  xor2s3
  U4110
  (
    .DIN1(n6467),
    .DIN1_t(n6467_t),
    .DIN2(n4846),
    .DIN2_t(n4846_t),
    .Q(n4845),
    .Q_t(n4845_t)
  );


  xor2s3
  U4111
  (
    .DIN1(n6465),
    .DIN1_t(n6465_t),
    .DIN2(n6466),
    .DIN2_t(n6466_t),
    .Q(n4846),
    .Q_t(n4846_t)
  );


  xor2s3
  U4112
  (
    .DIN1(n6552),
    .DIN1_t(n6552_t),
    .DIN2(n6710),
    .DIN2_t(n6710_t),
    .Q(n4844),
    .Q_t(n4844_t)
  );


  nnd2s3
  U4113
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2280),
    .DIN2_t(n2280_t),
    .Q(n4843),
    .Q_t(n4843_t)
  );


  xnr2s3
  U4114
  (
    .DIN1(n4847),
    .DIN1_t(n4847_t),
    .DIN2(n3095),
    .DIN2_t(n3095_t),
    .Q(DATA_9_6),
    .Q_t(DATA_9_6_t)
  );


  xnr2s3
  U4115
  (
    .DIN1(n4848),
    .DIN1_t(n4848_t),
    .DIN2(n4849),
    .DIN2_t(n4849_t),
    .Q(n3095),
    .Q_t(n3095_t)
  );


  xor2s3
  U4116
  (
    .DIN1(n6443),
    .DIN1_t(n6443_t),
    .DIN2(n4850),
    .DIN2_t(n4850_t),
    .Q(n4849),
    .Q_t(n4849_t)
  );


  xor2s3
  U4117
  (
    .DIN1(n6441),
    .DIN1_t(n6441_t),
    .DIN2(n6442),
    .DIN2_t(n6442_t),
    .Q(n4850),
    .Q_t(n4850_t)
  );


  xor2s3
  U4118
  (
    .DIN1(n6560),
    .DIN1_t(n6560_t),
    .DIN2(n6710),
    .DIN2_t(n6710_t),
    .Q(n4848),
    .Q_t(n4848_t)
  );


  nnd2s3
  U4119
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2279),
    .DIN2_t(n2279_t),
    .Q(n4847),
    .Q_t(n4847_t)
  );


  xnr2s3
  U4120
  (
    .DIN1(n4851),
    .DIN1_t(n4851_t),
    .DIN2(n3089),
    .DIN2_t(n3089_t),
    .Q(DATA_9_5),
    .Q_t(DATA_9_5_t)
  );


  xnr2s3
  U4121
  (
    .DIN1(n4852),
    .DIN1_t(n4852_t),
    .DIN2(n4853),
    .DIN2_t(n4853_t),
    .Q(n3089),
    .Q_t(n3089_t)
  );


  xor2s3
  U4122
  (
    .DIN1(n6461),
    .DIN1_t(n6461_t),
    .DIN2(n4854),
    .DIN2_t(n4854_t),
    .Q(n4853),
    .Q_t(n4853_t)
  );


  xor2s3
  U4123
  (
    .DIN1(n6459),
    .DIN1_t(n6459_t),
    .DIN2(n6460),
    .DIN2_t(n6460_t),
    .Q(n4854),
    .Q_t(n4854_t)
  );


  xor2s3
  U4124
  (
    .DIN1(n6554),
    .DIN1_t(n6554_t),
    .DIN2(n6709),
    .DIN2_t(n6709_t),
    .Q(n4852),
    .Q_t(n4852_t)
  );


  nnd2s3
  U4125
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2278),
    .DIN2_t(n2278_t),
    .Q(n4851),
    .Q_t(n4851_t)
  );


  xnr2s3
  U4126
  (
    .DIN1(n4855),
    .DIN1_t(n4855_t),
    .DIN2(n3083),
    .DIN2_t(n3083_t),
    .Q(DATA_9_4),
    .Q_t(DATA_9_4_t)
  );


  xnr2s3
  U4127
  (
    .DIN1(n4856),
    .DIN1_t(n4856_t),
    .DIN2(n4857),
    .DIN2_t(n4857_t),
    .Q(n3083),
    .Q_t(n3083_t)
  );


  xor2s3
  U4128
  (
    .DIN1(n6473),
    .DIN1_t(n6473_t),
    .DIN2(n4858),
    .DIN2_t(n4858_t),
    .Q(n4857),
    .Q_t(n4857_t)
  );


  xor2s3
  U4129
  (
    .DIN1(n6471),
    .DIN1_t(n6471_t),
    .DIN2(n6472),
    .DIN2_t(n6472_t),
    .Q(n4858),
    .Q_t(n4858_t)
  );


  xor2s3
  U4130
  (
    .DIN1(n6550),
    .DIN1_t(n6550_t),
    .DIN2(n6709),
    .DIN2_t(n6709_t),
    .Q(n4856),
    .Q_t(n4856_t)
  );


  nnd2s3
  U4131
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2277),
    .DIN2_t(n2277_t),
    .Q(n4855),
    .Q_t(n4855_t)
  );


  xnr2s3
  U4132
  (
    .DIN1(n4859),
    .DIN1_t(n4859_t),
    .DIN2(n3406),
    .DIN2_t(n3406_t),
    .Q(DATA_9_31),
    .Q_t(DATA_9_31_t)
  );


  xnr2s3
  U4133
  (
    .DIN1(n4860),
    .DIN1_t(n4860_t),
    .DIN2(n4861),
    .DIN2_t(n4861_t),
    .Q(n3406),
    .Q_t(n3406_t)
  );


  xor2s3
  U4134
  (
    .DIN1(n6533),
    .DIN1_t(n6533_t),
    .DIN2(n4862),
    .DIN2_t(n4862_t),
    .Q(n4861),
    .Q_t(n4861_t)
  );


  xor2s3
  U4135
  (
    .DIN1(n6531),
    .DIN1_t(n6531_t),
    .DIN2(n6532),
    .DIN2_t(n6532_t),
    .Q(n4862),
    .Q_t(n4862_t)
  );


  xor2s3
  U4136
  (
    .DIN1(n6534),
    .DIN1_t(n6534_t),
    .DIN2(n6696),
    .DIN2_t(n6696_t),
    .Q(n4860),
    .Q_t(n4860_t)
  );


  nnd2s3
  U4137
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2304),
    .DIN2_t(n2304_t),
    .Q(n4859),
    .Q_t(n4859_t)
  );


  xnr2s3
  U4138
  (
    .DIN1(n4863),
    .DIN1_t(n4863_t),
    .DIN2(n3388),
    .DIN2_t(n3388_t),
    .Q(DATA_9_30),
    .Q_t(DATA_9_30_t)
  );


  xnr2s3
  U4139
  (
    .DIN1(n4864),
    .DIN1_t(n4864_t),
    .DIN2(n4865),
    .DIN2_t(n4865_t),
    .Q(n3388),
    .Q_t(n3388_t)
  );


  xor2s3
  U4140
  (
    .DIN1(n6476),
    .DIN1_t(n6476_t),
    .DIN2(n4866),
    .DIN2_t(n4866_t),
    .Q(n4865),
    .Q_t(n4865_t)
  );


  xor2s3
  U4141
  (
    .DIN1(n6474),
    .DIN1_t(n6474_t),
    .DIN2(n6475),
    .DIN2_t(n6475_t),
    .Q(n4866),
    .Q_t(n4866_t)
  );


  xor2s3
  U4142
  (
    .DIN1(n6549),
    .DIN1_t(n6549_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4864),
    .Q_t(n4864_t)
  );


  nnd2s3
  U4143
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2303),
    .DIN2_t(n2303_t),
    .Q(n4863),
    .Q_t(n4863_t)
  );


  xnr2s3
  U4144
  (
    .DIN1(n4867),
    .DIN1_t(n4867_t),
    .DIN2(n3077),
    .DIN2_t(n3077_t),
    .Q(DATA_9_3),
    .Q_t(DATA_9_3_t)
  );


  xnr2s3
  U4145
  (
    .DIN1(n4868),
    .DIN1_t(n4868_t),
    .DIN2(n4869),
    .DIN2_t(n4869_t),
    .Q(n3077),
    .Q_t(n3077_t)
  );


  xor2s3
  U4146
  (
    .DIN1(n6470),
    .DIN1_t(n6470_t),
    .DIN2(n4870),
    .DIN2_t(n4870_t),
    .Q(n4869),
    .Q_t(n4869_t)
  );


  xor2s3
  U4147
  (
    .DIN1(n6468),
    .DIN1_t(n6468_t),
    .DIN2(n6469),
    .DIN2_t(n6469_t),
    .Q(n4870),
    .Q_t(n4870_t)
  );


  xor2s3
  U4148
  (
    .DIN1(n6551),
    .DIN1_t(n6551_t),
    .DIN2(n6709),
    .DIN2_t(n6709_t),
    .Q(n4868),
    .Q_t(n4868_t)
  );


  nnd2s3
  U4149
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2276),
    .DIN2_t(n2276_t),
    .Q(n4867),
    .Q_t(n4867_t)
  );


  xnr2s3
  U4150
  (
    .DIN1(n4871),
    .DIN1_t(n4871_t),
    .DIN2(n3371),
    .DIN2_t(n3371_t),
    .Q(DATA_9_29),
    .Q_t(DATA_9_29_t)
  );


  xnr2s3
  U4151
  (
    .DIN1(n4872),
    .DIN1_t(n4872_t),
    .DIN2(n4873),
    .DIN2_t(n4873_t),
    .Q(n3371),
    .Q_t(n3371_t)
  );


  xor2s3
  U4152
  (
    .DIN1(n6482),
    .DIN1_t(n6482_t),
    .DIN2(n4874),
    .DIN2_t(n4874_t),
    .Q(n4873),
    .Q_t(n4873_t)
  );


  xor2s3
  U4153
  (
    .DIN1(n6480),
    .DIN1_t(n6480_t),
    .DIN2(n6481),
    .DIN2_t(n6481_t),
    .Q(n4874),
    .Q_t(n4874_t)
  );


  xor2s3
  U4154
  (
    .DIN1(n6547),
    .DIN1_t(n6547_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4872),
    .Q_t(n4872_t)
  );


  nnd2s3
  U4155
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2302),
    .DIN2_t(n2302_t),
    .Q(n4871),
    .Q_t(n4871_t)
  );


  xnr2s3
  U4156
  (
    .DIN1(n4875),
    .DIN1_t(n4875_t),
    .DIN2(n3355),
    .DIN2_t(n3355_t),
    .Q(DATA_9_28),
    .Q_t(DATA_9_28_t)
  );


  xnr2s3
  U4157
  (
    .DIN1(n4876),
    .DIN1_t(n4876_t),
    .DIN2(n4877),
    .DIN2_t(n4877_t),
    .Q(n3355),
    .Q_t(n3355_t)
  );


  xor2s3
  U4158
  (
    .DIN1(n6485),
    .DIN1_t(n6485_t),
    .DIN2(n4878),
    .DIN2_t(n4878_t),
    .Q(n4877),
    .Q_t(n4877_t)
  );


  xor2s3
  U4159
  (
    .DIN1(n6483),
    .DIN1_t(n6483_t),
    .DIN2(n6484),
    .DIN2_t(n6484_t),
    .Q(n4878),
    .Q_t(n4878_t)
  );


  xor2s3
  U4160
  (
    .DIN1(n6546),
    .DIN1_t(n6546_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4876),
    .Q_t(n4876_t)
  );


  nnd2s3
  U4161
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2301),
    .DIN2_t(n2301_t),
    .Q(n4875),
    .Q_t(n4875_t)
  );


  xnr2s3
  U4162
  (
    .DIN1(n4879),
    .DIN1_t(n4879_t),
    .DIN2(n3349),
    .DIN2_t(n3349_t),
    .Q(DATA_9_27),
    .Q_t(DATA_9_27_t)
  );


  xnr2s3
  U4163
  (
    .DIN1(n4880),
    .DIN1_t(n4880_t),
    .DIN2(n4881),
    .DIN2_t(n4881_t),
    .Q(n3349),
    .Q_t(n3349_t)
  );


  xor2s3
  U4164
  (
    .DIN1(n6488),
    .DIN1_t(n6488_t),
    .DIN2(n4882),
    .DIN2_t(n4882_t),
    .Q(n4881),
    .Q_t(n4881_t)
  );


  xor2s3
  U4165
  (
    .DIN1(n6486),
    .DIN1_t(n6486_t),
    .DIN2(n6487),
    .DIN2_t(n6487_t),
    .Q(n4882),
    .Q_t(n4882_t)
  );


  xor2s3
  U4166
  (
    .DIN1(n6545),
    .DIN1_t(n6545_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4880),
    .Q_t(n4880_t)
  );


  nnd2s3
  U4167
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2300),
    .DIN2_t(n2300_t),
    .Q(n4879),
    .Q_t(n4879_t)
  );


  xnr2s3
  U4168
  (
    .DIN1(n4883),
    .DIN1_t(n4883_t),
    .DIN2(n3343),
    .DIN2_t(n3343_t),
    .Q(DATA_9_26),
    .Q_t(DATA_9_26_t)
  );


  xnr2s3
  U4169
  (
    .DIN1(n4884),
    .DIN1_t(n4884_t),
    .DIN2(n4885),
    .DIN2_t(n4885_t),
    .Q(n3343),
    .Q_t(n3343_t)
  );


  xor2s3
  U4170
  (
    .DIN1(n6494),
    .DIN1_t(n6494_t),
    .DIN2(n4886),
    .DIN2_t(n4886_t),
    .Q(n4885),
    .Q_t(n4885_t)
  );


  xor2s3
  U4171
  (
    .DIN1(n6492),
    .DIN1_t(n6492_t),
    .DIN2(n6493),
    .DIN2_t(n6493_t),
    .Q(n4886),
    .Q_t(n4886_t)
  );


  xor2s3
  U4172
  (
    .DIN1(n6543),
    .DIN1_t(n6543_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4884),
    .Q_t(n4884_t)
  );


  nnd2s3
  U4173
  (
    .DIN1(n6703),
    .DIN1_t(n6703_t),
    .DIN2(n2299),
    .DIN2_t(n2299_t),
    .Q(n4883),
    .Q_t(n4883_t)
  );


  xnr2s3
  U4174
  (
    .DIN1(n4887),
    .DIN1_t(n4887_t),
    .DIN2(n3337),
    .DIN2_t(n3337_t),
    .Q(DATA_9_25),
    .Q_t(DATA_9_25_t)
  );


  xnr2s3
  U4175
  (
    .DIN1(n4888),
    .DIN1_t(n4888_t),
    .DIN2(n4889),
    .DIN2_t(n4889_t),
    .Q(n3337),
    .Q_t(n3337_t)
  );


  xor2s3
  U4176
  (
    .DIN1(n6500),
    .DIN1_t(n6500_t),
    .DIN2(n4890),
    .DIN2_t(n4890_t),
    .Q(n4889),
    .Q_t(n4889_t)
  );


  xor2s3
  U4177
  (
    .DIN1(n6498),
    .DIN1_t(n6498_t),
    .DIN2(n6499),
    .DIN2_t(n6499_t),
    .Q(n4890),
    .Q_t(n4890_t)
  );


  xor2s3
  U4178
  (
    .DIN1(n6541),
    .DIN1_t(n6541_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4888),
    .Q_t(n4888_t)
  );


  nnd2s3
  U4179
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2298),
    .DIN2_t(n2298_t),
    .Q(n4887),
    .Q_t(n4887_t)
  );


  xnr2s3
  U4180
  (
    .DIN1(n4891),
    .DIN1_t(n4891_t),
    .DIN2(n3203),
    .DIN2_t(n3203_t),
    .Q(DATA_9_24),
    .Q_t(DATA_9_24_t)
  );


  xnr2s3
  U4181
  (
    .DIN1(n4892),
    .DIN1_t(n4892_t),
    .DIN2(n4893),
    .DIN2_t(n4893_t),
    .Q(n3203),
    .Q_t(n3203_t)
  );


  xor2s3
  U4182
  (
    .DIN1(n6503),
    .DIN1_t(n6503_t),
    .DIN2(n4894),
    .DIN2_t(n4894_t),
    .Q(n4893),
    .Q_t(n4893_t)
  );


  xor2s3
  U4183
  (
    .DIN1(n6501),
    .DIN1_t(n6501_t),
    .DIN2(n6502),
    .DIN2_t(n6502_t),
    .Q(n4894),
    .Q_t(n4894_t)
  );


  xor2s3
  U4184
  (
    .DIN1(n6540),
    .DIN1_t(n6540_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4892),
    .Q_t(n4892_t)
  );


  nnd2s3
  U4185
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2297),
    .DIN2_t(n2297_t),
    .Q(n4891),
    .Q_t(n4891_t)
  );


  xnr2s3
  U4186
  (
    .DIN1(n4895),
    .DIN1_t(n4895_t),
    .DIN2(n3197),
    .DIN2_t(n3197_t),
    .Q(DATA_9_23),
    .Q_t(DATA_9_23_t)
  );


  xnr2s3
  U4187
  (
    .DIN1(n4896),
    .DIN1_t(n4896_t),
    .DIN2(n4897),
    .DIN2_t(n4897_t),
    .Q(n3197),
    .Q_t(n3197_t)
  );


  xor2s3
  U4188
  (
    .DIN1(n6513),
    .DIN1_t(n6513_t),
    .DIN2(n4898),
    .DIN2_t(n4898_t),
    .Q(n4897),
    .Q_t(n4897_t)
  );


  xor2s3
  U4189
  (
    .DIN1(n6511),
    .DIN1_t(n6511_t),
    .DIN2(n6512),
    .DIN2_t(n6512_t),
    .Q(n4898),
    .Q_t(n4898_t)
  );


  xor2s3
  U4190
  (
    .DIN1(n6538),
    .DIN1_t(n6538_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4896),
    .Q_t(n4896_t)
  );


  nnd2s3
  U4191
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2296),
    .DIN2_t(n2296_t),
    .Q(n4895),
    .Q_t(n4895_t)
  );


  xnr2s3
  U4192
  (
    .DIN1(n4899),
    .DIN1_t(n4899_t),
    .DIN2(n3191),
    .DIN2_t(n3191_t),
    .Q(DATA_9_22),
    .Q_t(DATA_9_22_t)
  );


  xnr2s3
  U4193
  (
    .DIN1(n4900),
    .DIN1_t(n4900_t),
    .DIN2(n4901),
    .DIN2_t(n4901_t),
    .Q(n3191),
    .Q_t(n3191_t)
  );


  xor2s3
  U4194
  (
    .DIN1(n6516),
    .DIN1_t(n6516_t),
    .DIN2(n4902),
    .DIN2_t(n4902_t),
    .Q(n4901),
    .Q_t(n4901_t)
  );


  xor2s3
  U4195
  (
    .DIN1(n6514),
    .DIN1_t(n6514_t),
    .DIN2(n6515),
    .DIN2_t(n6515_t),
    .Q(n4902),
    .Q_t(n4902_t)
  );


  xor2s3
  U4196
  (
    .DIN1(n6537),
    .DIN1_t(n6537_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4900),
    .Q_t(n4900_t)
  );


  nnd2s3
  U4197
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2295),
    .DIN2_t(n2295_t),
    .Q(n4899),
    .Q_t(n4899_t)
  );


  xnr2s3
  U4198
  (
    .DIN1(n4903),
    .DIN1_t(n4903_t),
    .DIN2(n3185),
    .DIN2_t(n3185_t),
    .Q(DATA_9_21),
    .Q_t(DATA_9_21_t)
  );


  xnr2s3
  U4199
  (
    .DIN1(n4904),
    .DIN1_t(n4904_t),
    .DIN2(n4905),
    .DIN2_t(n4905_t),
    .Q(n3185),
    .Q_t(n3185_t)
  );


  xor2s3
  U4200
  (
    .DIN1(n6519),
    .DIN1_t(n6519_t),
    .DIN2(n4906),
    .DIN2_t(n4906_t),
    .Q(n4905),
    .Q_t(n4905_t)
  );


  xor2s3
  U4201
  (
    .DIN1(n6517),
    .DIN1_t(n6517_t),
    .DIN2(n6518),
    .DIN2_t(n6518_t),
    .Q(n4906),
    .Q_t(n4906_t)
  );


  xor2s3
  U4202
  (
    .DIN1(n6536),
    .DIN1_t(n6536_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4904),
    .Q_t(n4904_t)
  );


  nnd2s3
  U4203
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2294),
    .DIN2_t(n2294_t),
    .Q(n4903),
    .Q_t(n4903_t)
  );


  xnr2s3
  U4204
  (
    .DIN1(n4907),
    .DIN1_t(n4907_t),
    .DIN2(n3179),
    .DIN2_t(n3179_t),
    .Q(DATA_9_20),
    .Q_t(DATA_9_20_t)
  );


  xnr2s3
  U4205
  (
    .DIN1(n4908),
    .DIN1_t(n4908_t),
    .DIN2(n4909),
    .DIN2_t(n4909_t),
    .Q(n3179),
    .Q_t(n3179_t)
  );


  xor2s3
  U4206
  (
    .DIN1(n6522),
    .DIN1_t(n6522_t),
    .DIN2(n4910),
    .DIN2_t(n4910_t),
    .Q(n4909),
    .Q_t(n4909_t)
  );


  xor2s3
  U4207
  (
    .DIN1(n6520),
    .DIN1_t(n6520_t),
    .DIN2(n6521),
    .DIN2_t(n6521_t),
    .Q(n4910),
    .Q_t(n4910_t)
  );


  xor2s3
  U4208
  (
    .DIN1(n6535),
    .DIN1_t(n6535_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4908),
    .Q_t(n4908_t)
  );


  nnd2s3
  U4209
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2293),
    .DIN2_t(n2293_t),
    .Q(n4907),
    .Q_t(n4907_t)
  );


  xnr2s3
  U4210
  (
    .DIN1(n4911),
    .DIN1_t(n4911_t),
    .DIN2(n3071),
    .DIN2_t(n3071_t),
    .Q(DATA_9_2),
    .Q_t(DATA_9_2_t)
  );


  xnr2s3
  U4211
  (
    .DIN1(n4912),
    .DIN1_t(n4912_t),
    .DIN2(n4913),
    .DIN2_t(n4913_t),
    .Q(n3071),
    .Q_t(n3071_t)
  );


  xor2s3
  U4212
  (
    .DIN1(n6437),
    .DIN1_t(n6437_t),
    .DIN2(n4914),
    .DIN2_t(n4914_t),
    .Q(n4913),
    .Q_t(n4913_t)
  );


  xor2s3
  U4213
  (
    .DIN1(n6435),
    .DIN1_t(n6435_t),
    .DIN2(n6436),
    .DIN2_t(n6436_t),
    .Q(n4914),
    .Q_t(n4914_t)
  );


  xor2s3
  U4214
  (
    .DIN1(n6562),
    .DIN1_t(n6562_t),
    .DIN2(n6709),
    .DIN2_t(n6709_t),
    .Q(n4912),
    .Q_t(n4912_t)
  );


  nnd2s3
  U4215
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2275),
    .DIN2_t(n2275_t),
    .Q(n4911),
    .Q_t(n4911_t)
  );


  xnr2s3
  U4216
  (
    .DIN1(n4915),
    .DIN1_t(n4915_t),
    .DIN2(n3173),
    .DIN2_t(n3173_t),
    .Q(DATA_9_19),
    .Q_t(DATA_9_19_t)
  );


  xnr2s3
  U4217
  (
    .DIN1(n4916),
    .DIN1_t(n4916_t),
    .DIN2(n4917),
    .DIN2_t(n4917_t),
    .Q(n3173),
    .Q_t(n3173_t)
  );


  xor2s3
  U4218
  (
    .DIN1(n6479),
    .DIN1_t(n6479_t),
    .DIN2(n4918),
    .DIN2_t(n4918_t),
    .Q(n4917),
    .Q_t(n4917_t)
  );


  xor2s3
  U4219
  (
    .DIN1(n6477),
    .DIN1_t(n6477_t),
    .DIN2(n6478),
    .DIN2_t(n6478_t),
    .Q(n4918),
    .Q_t(n4918_t)
  );


  xor2s3
  U4220
  (
    .DIN1(n6548),
    .DIN1_t(n6548_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4916),
    .Q_t(n4916_t)
  );


  nnd2s3
  U4221
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2292),
    .DIN2_t(n2292_t),
    .Q(n4915),
    .Q_t(n4915_t)
  );


  xnr2s3
  U4222
  (
    .DIN1(n4919),
    .DIN1_t(n4919_t),
    .DIN2(n3167),
    .DIN2_t(n3167_t),
    .Q(DATA_9_18),
    .Q_t(DATA_9_18_t)
  );


  xnr2s3
  U4223
  (
    .DIN1(n4920),
    .DIN1_t(n4920_t),
    .DIN2(n4921),
    .DIN2_t(n4921_t),
    .Q(n3167),
    .Q_t(n3167_t)
  );


  xor2s3
  U4224
  (
    .DIN1(n6491),
    .DIN1_t(n6491_t),
    .DIN2(n4922),
    .DIN2_t(n4922_t),
    .Q(n4921),
    .Q_t(n4921_t)
  );


  xor2s3
  U4225
  (
    .DIN1(n6489),
    .DIN1_t(n6489_t),
    .DIN2(n6490),
    .DIN2_t(n6490_t),
    .Q(n4922),
    .Q_t(n4922_t)
  );


  xor2s3
  U4226
  (
    .DIN1(n6544),
    .DIN1_t(n6544_t),
    .DIN2(n6698),
    .DIN2_t(n6698_t),
    .Q(n4920),
    .Q_t(n4920_t)
  );


  nnd2s3
  U4227
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2291),
    .DIN2_t(n2291_t),
    .Q(n4919),
    .Q_t(n4919_t)
  );


  xnr2s3
  U4228
  (
    .DIN1(n4923),
    .DIN1_t(n4923_t),
    .DIN2(n3161),
    .DIN2_t(n3161_t),
    .Q(DATA_9_17),
    .Q_t(DATA_9_17_t)
  );


  xnr2s3
  U4229
  (
    .DIN1(n4924),
    .DIN1_t(n4924_t),
    .DIN2(n4925),
    .DIN2_t(n4925_t),
    .Q(n3161),
    .Q_t(n3161_t)
  );


  xor2s3
  U4230
  (
    .DIN1(n6497),
    .DIN1_t(n6497_t),
    .DIN2(n4926),
    .DIN2_t(n4926_t),
    .Q(n4925),
    .Q_t(n4925_t)
  );


  xor2s3
  U4231
  (
    .DIN1(n6495),
    .DIN1_t(n6495_t),
    .DIN2(n6496),
    .DIN2_t(n6496_t),
    .Q(n4926),
    .Q_t(n4926_t)
  );


  xor2s3
  U4232
  (
    .DIN1(n6542),
    .DIN1_t(n6542_t),
    .DIN2(n6697),
    .DIN2_t(n6697_t),
    .Q(n4924),
    .Q_t(n4924_t)
  );


  nnd2s3
  U4233
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2290),
    .DIN2_t(n2290_t),
    .Q(n4923),
    .Q_t(n4923_t)
  );


  xnr2s3
  U4234
  (
    .DIN1(n4927),
    .DIN1_t(n4927_t),
    .DIN2(n3155),
    .DIN2_t(n3155_t),
    .Q(DATA_9_16),
    .Q_t(DATA_9_16_t)
  );


  xnr2s3
  U4235
  (
    .DIN1(n4928),
    .DIN1_t(n4928_t),
    .DIN2(n4929),
    .DIN2_t(n4929_t),
    .Q(n3155),
    .Q_t(n3155_t)
  );


  xor2s3
  U4236
  (
    .DIN1(n6510),
    .DIN1_t(n6510_t),
    .DIN2(n4930),
    .DIN2_t(n4930_t),
    .Q(n4929),
    .Q_t(n4929_t)
  );


  xor2s3
  U4237
  (
    .DIN1(n6508),
    .DIN1_t(n6508_t),
    .DIN2(n6509),
    .DIN2_t(n6509_t),
    .Q(n4930),
    .Q_t(n4930_t)
  );


  xor2s3
  U4238
  (
    .DIN1(n6539),
    .DIN1_t(n6539_t),
    .DIN2(n6687),
    .DIN2_t(n6687_t),
    .Q(n4928),
    .Q_t(n4928_t)
  );


  nnd2s3
  U4239
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2289),
    .DIN2_t(n2289_t),
    .Q(n4927),
    .Q_t(n4927_t)
  );


  xnr2s3
  U4240
  (
    .DIN1(n4931),
    .DIN1_t(n4931_t),
    .DIN2(n3149),
    .DIN2_t(n3149_t),
    .Q(DATA_9_15),
    .Q_t(DATA_9_15_t)
  );


  xnr2s3
  U4241
  (
    .DIN1(n4932),
    .DIN1_t(n4932_t),
    .DIN2(n4933),
    .DIN2_t(n4933_t),
    .Q(n3149),
    .Q_t(n3149_t)
  );


  xor2s3
  U4242
  (
    .DIN1(n6440),
    .DIN1_t(n6440_t),
    .DIN2(n4934),
    .DIN2_t(n4934_t),
    .Q(n4933),
    .Q_t(n4933_t)
  );


  xor2s3
  U4243
  (
    .DIN1(n6438),
    .DIN1_t(n6438_t),
    .DIN2(n6439),
    .DIN2_t(n6439_t),
    .Q(n4934),
    .Q_t(n4934_t)
  );


  xor2s3
  U4244
  (
    .DIN1(n6561),
    .DIN1_t(n6561_t),
    .DIN2(n6708),
    .DIN2_t(n6708_t),
    .Q(n4932),
    .Q_t(n4932_t)
  );


  nnd2s3
  U4245
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2288),
    .DIN2_t(n2288_t),
    .Q(n4931),
    .Q_t(n4931_t)
  );


  xnr2s3
  U4246
  (
    .DIN1(n4935),
    .DIN1_t(n4935_t),
    .DIN2(n3143),
    .DIN2_t(n3143_t),
    .Q(DATA_9_14),
    .Q_t(DATA_9_14_t)
  );


  xnr2s3
  U4247
  (
    .DIN1(n4936),
    .DIN1_t(n4936_t),
    .DIN2(n4937),
    .DIN2_t(n4937_t),
    .Q(n3143),
    .Q_t(n3143_t)
  );


  xor2s3
  U4248
  (
    .DIN1(n6525),
    .DIN1_t(n6525_t),
    .DIN2(n4938),
    .DIN2_t(n4938_t),
    .Q(n4937),
    .Q_t(n4937_t)
  );


  xor2s3
  U4249
  (
    .DIN1(n6523),
    .DIN1_t(n6523_t),
    .DIN2(n6524),
    .DIN2_t(n6524_t),
    .Q(n4938),
    .Q_t(n4938_t)
  );


  xor2s3
  U4250
  (
    .DIN1(n6526),
    .DIN1_t(n6526_t),
    .DIN2(n6708),
    .DIN2_t(n6708_t),
    .Q(n4936),
    .Q_t(n4936_t)
  );


  nnd2s3
  U4251
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2287),
    .DIN2_t(n2287_t),
    .Q(n4935),
    .Q_t(n4935_t)
  );


  xnr2s3
  U4252
  (
    .DIN1(n4939),
    .DIN1_t(n4939_t),
    .DIN2(n3137),
    .DIN2_t(n3137_t),
    .Q(DATA_9_13),
    .Q_t(DATA_9_13_t)
  );


  xnr2s3
  U4253
  (
    .DIN1(n4940),
    .DIN1_t(n4940_t),
    .DIN2(n4941),
    .DIN2_t(n4941_t),
    .Q(n3137),
    .Q_t(n3137_t)
  );


  xor2s3
  U4254
  (
    .DIN1(n6449),
    .DIN1_t(n6449_t),
    .DIN2(n4942),
    .DIN2_t(n4942_t),
    .Q(n4941),
    .Q_t(n4941_t)
  );


  xor2s3
  U4255
  (
    .DIN1(n6447),
    .DIN1_t(n6447_t),
    .DIN2(n6448),
    .DIN2_t(n6448_t),
    .Q(n4942),
    .Q_t(n4942_t)
  );


  xor2s3
  U4256
  (
    .DIN1(n6558),
    .DIN1_t(n6558_t),
    .DIN2(n6708),
    .DIN2_t(n6708_t),
    .Q(n4940),
    .Q_t(n4940_t)
  );


  nnd2s3
  U4257
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2286),
    .DIN2_t(n2286_t),
    .Q(n4939),
    .Q_t(n4939_t)
  );


  xnr2s3
  U4258
  (
    .DIN1(n4943),
    .DIN1_t(n4943_t),
    .DIN2(n3131),
    .DIN2_t(n3131_t),
    .Q(DATA_9_12),
    .Q_t(DATA_9_12_t)
  );


  xnr2s3
  U4259
  (
    .DIN1(n4944),
    .DIN1_t(n4944_t),
    .DIN2(n4945),
    .DIN2_t(n4945_t),
    .Q(n3131),
    .Q_t(n3131_t)
  );


  xor2s3
  U4260
  (
    .DIN1(n6458),
    .DIN1_t(n6458_t),
    .DIN2(n4946),
    .DIN2_t(n4946_t),
    .Q(n4945),
    .Q_t(n4945_t)
  );


  xor2s3
  U4261
  (
    .DIN1(n6456),
    .DIN1_t(n6456_t),
    .DIN2(n6457),
    .DIN2_t(n6457_t),
    .Q(n4946),
    .Q_t(n4946_t)
  );


  xor2s3
  U4262
  (
    .DIN1(n6555),
    .DIN1_t(n6555_t),
    .DIN2(n6708),
    .DIN2_t(n6708_t),
    .Q(n4944),
    .Q_t(n4944_t)
  );


  nnd2s3
  U4263
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2285),
    .DIN2_t(n2285_t),
    .Q(n4943),
    .Q_t(n4943_t)
  );


  xnr2s3
  U4264
  (
    .DIN1(n4947),
    .DIN1_t(n4947_t),
    .DIN2(n3125),
    .DIN2_t(n3125_t),
    .Q(DATA_9_11),
    .Q_t(DATA_9_11_t)
  );


  xnr2s3
  U4265
  (
    .DIN1(n4948),
    .DIN1_t(n4948_t),
    .DIN2(n4949),
    .DIN2_t(n4949_t),
    .Q(n3125),
    .Q_t(n3125_t)
  );


  xor2s3
  U4266
  (
    .DIN1(n6446),
    .DIN1_t(n6446_t),
    .DIN2(n4950),
    .DIN2_t(n4950_t),
    .Q(n4949),
    .Q_t(n4949_t)
  );


  xor2s3
  U4267
  (
    .DIN1(n6444),
    .DIN1_t(n6444_t),
    .DIN2(n6445),
    .DIN2_t(n6445_t),
    .Q(n4950),
    .Q_t(n4950_t)
  );


  xor2s3
  U4268
  (
    .DIN1(n6559),
    .DIN1_t(n6559_t),
    .DIN2(n6707),
    .DIN2_t(n6707_t),
    .Q(n4948),
    .Q_t(n4948_t)
  );


  nnd2s3
  U4269
  (
    .DIN1(n6704),
    .DIN1_t(n6704_t),
    .DIN2(n2284),
    .DIN2_t(n2284_t),
    .Q(n4947),
    .Q_t(n4947_t)
  );


  xnr2s3
  U4270
  (
    .DIN1(n4951),
    .DIN1_t(n4951_t),
    .DIN2(n3119),
    .DIN2_t(n3119_t),
    .Q(DATA_9_10),
    .Q_t(DATA_9_10_t)
  );


  xnr2s3
  U4271
  (
    .DIN1(n4952),
    .DIN1_t(n4952_t),
    .DIN2(n4953),
    .DIN2_t(n4953_t),
    .Q(n3119),
    .Q_t(n3119_t)
  );


  xor2s3
  U4272
  (
    .DIN1(n6452),
    .DIN1_t(n6452_t),
    .DIN2(n4954),
    .DIN2_t(n4954_t),
    .Q(n4953),
    .Q_t(n4953_t)
  );


  xor2s3
  U4273
  (
    .DIN1(n6450),
    .DIN1_t(n6450_t),
    .DIN2(n6451),
    .DIN2_t(n6451_t),
    .Q(n4954),
    .Q_t(n4954_t)
  );


  xor2s3
  U4274
  (
    .DIN1(n6557),
    .DIN1_t(n6557_t),
    .DIN2(n6707),
    .DIN2_t(n6707_t),
    .Q(n4952),
    .Q_t(n4952_t)
  );


  nnd2s3
  U4275
  (
    .DIN1(n6705),
    .DIN1_t(n6705_t),
    .DIN2(n2283),
    .DIN2_t(n2283_t),
    .Q(n4951),
    .Q_t(n4951_t)
  );


  xnr2s3
  U4276
  (
    .DIN1(n4955),
    .DIN1_t(n4955_t),
    .DIN2(n3065),
    .DIN2_t(n3065_t),
    .Q(DATA_9_1),
    .Q_t(DATA_9_1_t)
  );


  xnr2s3
  U4277
  (
    .DIN1(n4956),
    .DIN1_t(n4956_t),
    .DIN2(n4957),
    .DIN2_t(n4957_t),
    .Q(n3065),
    .Q_t(n3065_t)
  );


  xor2s3
  U4278
  (
    .DIN1(n6529),
    .DIN1_t(n6529_t),
    .DIN2(n4958),
    .DIN2_t(n4958_t),
    .Q(n4957),
    .Q_t(n4957_t)
  );


  xor2s3
  U4279
  (
    .DIN1(n6527),
    .DIN1_t(n6527_t),
    .DIN2(n6528),
    .DIN2_t(n6528_t),
    .Q(n4958),
    .Q_t(n4958_t)
  );


  xor2s3
  U4280
  (
    .DIN1(n6530),
    .DIN1_t(n6530_t),
    .DIN2(n6707),
    .DIN2_t(n6707_t),
    .Q(n4956),
    .Q_t(n4956_t)
  );


  nnd2s3
  U4281
  (
    .DIN1(n6705),
    .DIN1_t(n6705_t),
    .DIN2(n2274),
    .DIN2_t(n2274_t),
    .Q(n4955),
    .Q_t(n4955_t)
  );


  xnr2s3
  U4282
  (
    .DIN1(n4959),
    .DIN1_t(n4959_t),
    .DIN2(n3059),
    .DIN2_t(n3059_t),
    .Q(DATA_9_0),
    .Q_t(DATA_9_0_t)
  );


  xnr2s3
  U4283
  (
    .DIN1(n4960),
    .DIN1_t(n4960_t),
    .DIN2(n4961),
    .DIN2_t(n4961_t),
    .Q(n3059),
    .Q_t(n3059_t)
  );


  xor2s3
  U4284
  (
    .DIN1(n6464),
    .DIN1_t(n6464_t),
    .DIN2(n4962),
    .DIN2_t(n4962_t),
    .Q(n4961),
    .Q_t(n4961_t)
  );


  xor2s3
  U4285
  (
    .DIN1(n6462),
    .DIN1_t(n6462_t),
    .DIN2(n6463),
    .DIN2_t(n6463_t),
    .Q(n4962),
    .Q_t(n4962_t)
  );


  xor2s3
  U4286
  (
    .DIN1(n6553),
    .DIN1_t(n6553_t),
    .DIN2(n6707),
    .DIN2_t(n6707_t),
    .Q(n4960),
    .Q_t(n4960_t)
  );


  nnd2s3
  U4287
  (
    .DIN1(n6705),
    .DIN1_t(n6705_t),
    .DIN2(n2273),
    .DIN2_t(n2273_t),
    .Q(n4959),
    .Q_t(n4959_t)
  );


  i1s3
  U4288
  (
    .DIN(n6337),
    .DIN_t(n6337_t),
    .Q(n1729),
    .Q_t(n1729_t)
  );


  i1s3
  U4289
  (
    .DIN(n6336),
    .DIN_t(n6336_t),
    .Q(n1730),
    .Q_t(n1730_t)
  );


  i1s3
  U4290
  (
    .DIN(n6331),
    .DIN_t(n6331_t),
    .Q(n1731),
    .Q_t(n1731_t)
  );


  i1s3
  U4291
  (
    .DIN(n6326),
    .DIN_t(n6326_t),
    .Q(n1732),
    .Q_t(n1732_t)
  );


  i1s3
  U4292
  (
    .DIN(n6321),
    .DIN_t(n6321_t),
    .Q(n1733),
    .Q_t(n1733_t)
  );


  i1s3
  U4293
  (
    .DIN(n6316),
    .DIN_t(n6316_t),
    .Q(n1734),
    .Q_t(n1734_t)
  );


  i1s3
  U4294
  (
    .DIN(n6311),
    .DIN_t(n6311_t),
    .Q(n1735),
    .Q_t(n1735_t)
  );


  i1s3
  U4295
  (
    .DIN(n6306),
    .DIN_t(n6306_t),
    .Q(n1736),
    .Q_t(n1736_t)
  );


  i1s3
  U4296
  (
    .DIN(n6301),
    .DIN_t(n6301_t),
    .Q(n1737),
    .Q_t(n1737_t)
  );


  i1s3
  U4297
  (
    .DIN(n6296),
    .DIN_t(n6296_t),
    .Q(n1738),
    .Q_t(n1738_t)
  );


  i1s3
  U4298
  (
    .DIN(n6291),
    .DIN_t(n6291_t),
    .Q(n1739),
    .Q_t(n1739_t)
  );


  i1s3
  U4299
  (
    .DIN(n6285),
    .DIN_t(n6285_t),
    .Q(n1740),
    .Q_t(n1740_t)
  );


  i1s3
  U4300
  (
    .DIN(n6280),
    .DIN_t(n6280_t),
    .Q(n1741),
    .Q_t(n1741_t)
  );


  i1s3
  U4301
  (
    .DIN(n6275),
    .DIN_t(n6275_t),
    .Q(n1742),
    .Q_t(n1742_t)
  );


  i1s3
  U4302
  (
    .DIN(n6270),
    .DIN_t(n6270_t),
    .Q(n1743),
    .Q_t(n1743_t)
  );


  i1s3
  U4303
  (
    .DIN(n6265),
    .DIN_t(n6265_t),
    .Q(n1744),
    .Q_t(n1744_t)
  );


  i1s3
  U4304
  (
    .DIN(n6260),
    .DIN_t(n6260_t),
    .Q(n1745),
    .Q_t(n1745_t)
  );


  i1s3
  U4305
  (
    .DIN(n6256),
    .DIN_t(n6256_t),
    .Q(n1746),
    .Q_t(n1746_t)
  );


  i1s3
  U4306
  (
    .DIN(n6252),
    .DIN_t(n6252_t),
    .Q(n1747),
    .Q_t(n1747_t)
  );


  i1s3
  U4307
  (
    .DIN(n6248),
    .DIN_t(n6248_t),
    .Q(n1748),
    .Q_t(n1748_t)
  );


  i1s3
  U4308
  (
    .DIN(n6244),
    .DIN_t(n6244_t),
    .Q(n1749),
    .Q_t(n1749_t)
  );


  i1s3
  U4309
  (
    .DIN(n6240),
    .DIN_t(n6240_t),
    .Q(n1750),
    .Q_t(n1750_t)
  );


  i1s3
  U4310
  (
    .DIN(n6236),
    .DIN_t(n6236_t),
    .Q(n1751),
    .Q_t(n1751_t)
  );


  i1s3
  U4311
  (
    .DIN(n6232),
    .DIN_t(n6232_t),
    .Q(n1752),
    .Q_t(n1752_t)
  );


  i1s3
  U4312
  (
    .DIN(n6228),
    .DIN_t(n6228_t),
    .Q(n1753),
    .Q_t(n1753_t)
  );


  i1s3
  U4313
  (
    .DIN(n6224),
    .DIN_t(n6224_t),
    .Q(n1754),
    .Q_t(n1754_t)
  );


  i1s3
  U4314
  (
    .DIN(n6220),
    .DIN_t(n6220_t),
    .Q(n1755),
    .Q_t(n1755_t)
  );


  i1s3
  U4315
  (
    .DIN(n6216),
    .DIN_t(n6216_t),
    .Q(n1756),
    .Q_t(n1756_t)
  );


  i1s3
  U4316
  (
    .DIN(n6212),
    .DIN_t(n6212_t),
    .Q(n1757),
    .Q_t(n1757_t)
  );


  i1s3
  U4317
  (
    .DIN(n6208),
    .DIN_t(n6208_t),
    .Q(n1758),
    .Q_t(n1758_t)
  );


  i1s3
  U4318
  (
    .DIN(n6204),
    .DIN_t(n6204_t),
    .Q(n1759),
    .Q_t(n1759_t)
  );


  i1s3
  U4319
  (
    .DIN(n6200),
    .DIN_t(n6200_t),
    .Q(n1760),
    .Q_t(n1760_t)
  );


  i1s3
  U4320
  (
    .DIN(n6344),
    .DIN_t(n6344_t),
    .Q(n1761),
    .Q_t(n1761_t)
  );


  i1s3
  U4321
  (
    .DIN(n6345),
    .DIN_t(n6345_t),
    .Q(n1762),
    .Q_t(n1762_t)
  );


  i1s3
  U4322
  (
    .DIN(n6346),
    .DIN_t(n6346_t),
    .Q(n1763),
    .Q_t(n1763_t)
  );


  i1s3
  U4323
  (
    .DIN(n6347),
    .DIN_t(n6347_t),
    .Q(n1764),
    .Q_t(n1764_t)
  );


  i1s3
  U4324
  (
    .DIN(n6348),
    .DIN_t(n6348_t),
    .Q(n1765),
    .Q_t(n1765_t)
  );


  i1s3
  U4325
  (
    .DIN(n6349),
    .DIN_t(n6349_t),
    .Q(n1766),
    .Q_t(n1766_t)
  );


  i1s3
  U4326
  (
    .DIN(n6350),
    .DIN_t(n6350_t),
    .Q(n1767),
    .Q_t(n1767_t)
  );


  i1s3
  U4327
  (
    .DIN(n6351),
    .DIN_t(n6351_t),
    .Q(n1768),
    .Q_t(n1768_t)
  );


  i1s3
  U4328
  (
    .DIN(n6352),
    .DIN_t(n6352_t),
    .Q(n1769),
    .Q_t(n1769_t)
  );


  i1s3
  U4329
  (
    .DIN(n6353),
    .DIN_t(n6353_t),
    .Q(n1770),
    .Q_t(n1770_t)
  );


  i1s3
  U4330
  (
    .DIN(n6355),
    .DIN_t(n6355_t),
    .Q(n1771),
    .Q_t(n1771_t)
  );


  i1s3
  U4331
  (
    .DIN(n6356),
    .DIN_t(n6356_t),
    .Q(n1772),
    .Q_t(n1772_t)
  );


  i1s3
  U4332
  (
    .DIN(n6357),
    .DIN_t(n6357_t),
    .Q(n1773),
    .Q_t(n1773_t)
  );


  i1s3
  U4333
  (
    .DIN(n6358),
    .DIN_t(n6358_t),
    .Q(n1774),
    .Q_t(n1774_t)
  );


  i1s3
  U4334
  (
    .DIN(n6359),
    .DIN_t(n6359_t),
    .Q(n1775),
    .Q_t(n1775_t)
  );


  i1s3
  U4335
  (
    .DIN(n6360),
    .DIN_t(n6360_t),
    .Q(n1776),
    .Q_t(n1776_t)
  );


  i1s3
  U4336
  (
    .DIN(n6361),
    .DIN_t(n6361_t),
    .Q(n1777),
    .Q_t(n1777_t)
  );


  i1s3
  U4337
  (
    .DIN(n6362),
    .DIN_t(n6362_t),
    .Q(n1778),
    .Q_t(n1778_t)
  );


  i1s3
  U4338
  (
    .DIN(n6363),
    .DIN_t(n6363_t),
    .Q(n1779),
    .Q_t(n1779_t)
  );


  i1s3
  U4339
  (
    .DIN(n6364),
    .DIN_t(n6364_t),
    .Q(n1780),
    .Q_t(n1780_t)
  );


  i1s3
  U4340
  (
    .DIN(n6365),
    .DIN_t(n6365_t),
    .Q(n1781),
    .Q_t(n1781_t)
  );


  i1s3
  U4341
  (
    .DIN(n6366),
    .DIN_t(n6366_t),
    .Q(n1782),
    .Q_t(n1782_t)
  );


  i1s3
  U4342
  (
    .DIN(n6367),
    .DIN_t(n6367_t),
    .Q(n1783),
    .Q_t(n1783_t)
  );


  i1s3
  U4343
  (
    .DIN(n6368),
    .DIN_t(n6368_t),
    .Q(n1784),
    .Q_t(n1784_t)
  );


  i1s3
  U4344
  (
    .DIN(n6369),
    .DIN_t(n6369_t),
    .Q(n1785),
    .Q_t(n1785_t)
  );


  i1s3
  U4345
  (
    .DIN(n6370),
    .DIN_t(n6370_t),
    .Q(n1786),
    .Q_t(n1786_t)
  );


  i1s3
  U4346
  (
    .DIN(n6371),
    .DIN_t(n6371_t),
    .Q(n1787),
    .Q_t(n1787_t)
  );


  i1s3
  U4347
  (
    .DIN(n6372),
    .DIN_t(n6372_t),
    .Q(n1788),
    .Q_t(n1788_t)
  );


  i1s3
  U4348
  (
    .DIN(n6373),
    .DIN_t(n6373_t),
    .Q(n1789),
    .Q_t(n1789_t)
  );


  i1s3
  U4349
  (
    .DIN(n6374),
    .DIN_t(n6374_t),
    .Q(n1790),
    .Q_t(n1790_t)
  );


  i1s3
  U4350
  (
    .DIN(n6375),
    .DIN_t(n6375_t),
    .Q(n1791),
    .Q_t(n1791_t)
  );


  i1s3
  U4351
  (
    .DIN(n6343),
    .DIN_t(n6343_t),
    .Q(n1792),
    .Q_t(n1792_t)
  );


  i1s3
  U4352
  (
    .DIN(n6430),
    .DIN_t(n6430_t),
    .Q(n1793),
    .Q_t(n1793_t)
  );


  i1s3
  U4353
  (
    .DIN(n6383),
    .DIN_t(n6383_t),
    .Q(n1794),
    .Q_t(n1794_t)
  );


  i1s3
  U4354
  (
    .DIN(n6385),
    .DIN_t(n6385_t),
    .Q(n1795),
    .Q_t(n1795_t)
  );


  i1s3
  U4355
  (
    .DIN(n6387),
    .DIN_t(n6387_t),
    .Q(n1796),
    .Q_t(n1796_t)
  );


  i1s3
  U4356
  (
    .DIN(n6389),
    .DIN_t(n6389_t),
    .Q(n1797),
    .Q_t(n1797_t)
  );


  i1s3
  U4357
  (
    .DIN(n6391),
    .DIN_t(n6391_t),
    .Q(n1798),
    .Q_t(n1798_t)
  );


  i1s3
  U4358
  (
    .DIN(n6393),
    .DIN_t(n6393_t),
    .Q(n1799),
    .Q_t(n1799_t)
  );


  i1s3
  U4359
  (
    .DIN(n6395),
    .DIN_t(n6395_t),
    .Q(n1800),
    .Q_t(n1800_t)
  );


  i1s3
  U4360
  (
    .DIN(n6397),
    .DIN_t(n6397_t),
    .Q(n1801),
    .Q_t(n1801_t)
  );


  i1s3
  U4361
  (
    .DIN(n6399),
    .DIN_t(n6399_t),
    .Q(n1802),
    .Q_t(n1802_t)
  );


  i1s3
  U4362
  (
    .DIN(n6401),
    .DIN_t(n6401_t),
    .Q(n1803),
    .Q_t(n1803_t)
  );


  i1s3
  U4363
  (
    .DIN(n6403),
    .DIN_t(n6403_t),
    .Q(n1804),
    .Q_t(n1804_t)
  );


  i1s3
  U4364
  (
    .DIN(n6405),
    .DIN_t(n6405_t),
    .Q(n1805),
    .Q_t(n1805_t)
  );


  i1s3
  U4365
  (
    .DIN(n6407),
    .DIN_t(n6407_t),
    .Q(n1806),
    .Q_t(n1806_t)
  );


  i1s3
  U4366
  (
    .DIN(n6409),
    .DIN_t(n6409_t),
    .Q(n1807),
    .Q_t(n1807_t)
  );


  i1s3
  U4367
  (
    .DIN(n6411),
    .DIN_t(n6411_t),
    .Q(n1808),
    .Q_t(n1808_t)
  );


  i1s3
  U4368
  (
    .DIN(n6413),
    .DIN_t(n6413_t),
    .Q(n1809),
    .Q_t(n1809_t)
  );


  i1s3
  U4369
  (
    .DIN(n6415),
    .DIN_t(n6415_t),
    .Q(n1810),
    .Q_t(n1810_t)
  );


  i1s3
  U4370
  (
    .DIN(n6416),
    .DIN_t(n6416_t),
    .Q(n1811),
    .Q_t(n1811_t)
  );


  i1s3
  U4371
  (
    .DIN(n6417),
    .DIN_t(n6417_t),
    .Q(n1812),
    .Q_t(n1812_t)
  );


  i1s3
  U4372
  (
    .DIN(n6418),
    .DIN_t(n6418_t),
    .Q(n1813),
    .Q_t(n1813_t)
  );


  i1s3
  U4373
  (
    .DIN(n6419),
    .DIN_t(n6419_t),
    .Q(n1814),
    .Q_t(n1814_t)
  );


  i1s3
  U4374
  (
    .DIN(n6420),
    .DIN_t(n6420_t),
    .Q(n1815),
    .Q_t(n1815_t)
  );


  i1s3
  U4375
  (
    .DIN(n6421),
    .DIN_t(n6421_t),
    .Q(n1816),
    .Q_t(n1816_t)
  );


  i1s3
  U4376
  (
    .DIN(n6422),
    .DIN_t(n6422_t),
    .Q(n1817),
    .Q_t(n1817_t)
  );


  i1s3
  U4377
  (
    .DIN(n6423),
    .DIN_t(n6423_t),
    .Q(n1818),
    .Q_t(n1818_t)
  );


  i1s3
  U4378
  (
    .DIN(n6424),
    .DIN_t(n6424_t),
    .Q(n1819),
    .Q_t(n1819_t)
  );


  i1s3
  U4379
  (
    .DIN(n6425),
    .DIN_t(n6425_t),
    .Q(n1820),
    .Q_t(n1820_t)
  );


  i1s3
  U4380
  (
    .DIN(n6426),
    .DIN_t(n6426_t),
    .Q(n1821),
    .Q_t(n1821_t)
  );


  i1s3
  U4381
  (
    .DIN(n6427),
    .DIN_t(n6427_t),
    .Q(n1822),
    .Q_t(n1822_t)
  );


  i1s3
  U4382
  (
    .DIN(n6428),
    .DIN_t(n6428_t),
    .Q(n1823),
    .Q_t(n1823_t)
  );


  i1s3
  U4383
  (
    .DIN(n6429),
    .DIN_t(n6429_t),
    .Q(n1824),
    .Q_t(n1824_t)
  );


  i1s3
  U4384
  (
    .DIN(n4964),
    .DIN_t(n4964_t),
    .Q(n1825),
    .Q_t(n1825_t)
  );


  i1s3
  U4385
  (
    .DIN(n4965),
    .DIN_t(n4965_t),
    .Q(n1826),
    .Q_t(n1826_t)
  );


  i1s3
  U4386
  (
    .DIN(n4966),
    .DIN_t(n4966_t),
    .Q(n1827),
    .Q_t(n1827_t)
  );


  i1s3
  U4387
  (
    .DIN(n4967),
    .DIN_t(n4967_t),
    .Q(n1828),
    .Q_t(n1828_t)
  );


  i1s3
  U4388
  (
    .DIN(n4968),
    .DIN_t(n4968_t),
    .Q(n1829),
    .Q_t(n1829_t)
  );


  i1s3
  U4389
  (
    .DIN(n4969),
    .DIN_t(n4969_t),
    .Q(n1830),
    .Q_t(n1830_t)
  );


  i1s3
  U4390
  (
    .DIN(n4970),
    .DIN_t(n4970_t),
    .Q(n1831),
    .Q_t(n1831_t)
  );


  i1s3
  U4391
  (
    .DIN(n4971),
    .DIN_t(n4971_t),
    .Q(n1832),
    .Q_t(n1832_t)
  );


  i1s3
  U4392
  (
    .DIN(n4972),
    .DIN_t(n4972_t),
    .Q(n1833),
    .Q_t(n1833_t)
  );


  i1s3
  U4393
  (
    .DIN(n4973),
    .DIN_t(n4973_t),
    .Q(n1834),
    .Q_t(n1834_t)
  );


  i1s3
  U4394
  (
    .DIN(n4974),
    .DIN_t(n4974_t),
    .Q(n1835),
    .Q_t(n1835_t)
  );


  i1s3
  U4395
  (
    .DIN(n4975),
    .DIN_t(n4975_t),
    .Q(n1836),
    .Q_t(n1836_t)
  );


  i1s3
  U4396
  (
    .DIN(n4976),
    .DIN_t(n4976_t),
    .Q(n1837),
    .Q_t(n1837_t)
  );


  i1s3
  U4397
  (
    .DIN(n4977),
    .DIN_t(n4977_t),
    .Q(n1838),
    .Q_t(n1838_t)
  );


  i1s3
  U4398
  (
    .DIN(n4978),
    .DIN_t(n4978_t),
    .Q(n1839),
    .Q_t(n1839_t)
  );


  i1s3
  U4399
  (
    .DIN(n4979),
    .DIN_t(n4979_t),
    .Q(n1840),
    .Q_t(n1840_t)
  );


  i1s3
  U4400
  (
    .DIN(n4980),
    .DIN_t(n4980_t),
    .Q(n1841),
    .Q_t(n1841_t)
  );


  i1s3
  U4401
  (
    .DIN(n4981),
    .DIN_t(n4981_t),
    .Q(n1842),
    .Q_t(n1842_t)
  );


  i1s3
  U4402
  (
    .DIN(n4982),
    .DIN_t(n4982_t),
    .Q(n1843),
    .Q_t(n1843_t)
  );


  i1s3
  U4403
  (
    .DIN(n4983),
    .DIN_t(n4983_t),
    .Q(n1844),
    .Q_t(n1844_t)
  );


  i1s3
  U4404
  (
    .DIN(n4984),
    .DIN_t(n4984_t),
    .Q(n1845),
    .Q_t(n1845_t)
  );


  i1s3
  U4405
  (
    .DIN(n4985),
    .DIN_t(n4985_t),
    .Q(n1846),
    .Q_t(n1846_t)
  );


  i1s3
  U4406
  (
    .DIN(n4986),
    .DIN_t(n4986_t),
    .Q(n1847),
    .Q_t(n1847_t)
  );


  i1s3
  U4407
  (
    .DIN(n4987),
    .DIN_t(n4987_t),
    .Q(n1848),
    .Q_t(n1848_t)
  );


  i1s3
  U4408
  (
    .DIN(n4988),
    .DIN_t(n4988_t),
    .Q(n1849),
    .Q_t(n1849_t)
  );


  i1s3
  U4409
  (
    .DIN(n4989),
    .DIN_t(n4989_t),
    .Q(n1850),
    .Q_t(n1850_t)
  );


  i1s3
  U4410
  (
    .DIN(n4990),
    .DIN_t(n4990_t),
    .Q(n1851),
    .Q_t(n1851_t)
  );


  i1s3
  U4411
  (
    .DIN(n4991),
    .DIN_t(n4991_t),
    .Q(n1852),
    .Q_t(n1852_t)
  );


  i1s3
  U4412
  (
    .DIN(n4992),
    .DIN_t(n4992_t),
    .Q(n1853),
    .Q_t(n1853_t)
  );


  i1s3
  U4413
  (
    .DIN(n4993),
    .DIN_t(n4993_t),
    .Q(n1854),
    .Q_t(n1854_t)
  );


  i1s3
  U4414
  (
    .DIN(n4994),
    .DIN_t(n4994_t),
    .Q(n1855),
    .Q_t(n1855_t)
  );


  i1s3
  U4415
  (
    .DIN(n4963),
    .DIN_t(n4963_t),
    .Q(n1856),
    .Q_t(n1856_t)
  );


  i1s3
  U4416
  (
    .DIN(n5122),
    .DIN_t(n5122_t),
    .Q(n1857),
    .Q_t(n1857_t)
  );


  i1s3
  U4417
  (
    .DIN(n5118),
    .DIN_t(n5118_t),
    .Q(n1858),
    .Q_t(n1858_t)
  );


  i1s3
  U4418
  (
    .DIN(n5114),
    .DIN_t(n5114_t),
    .Q(n1859),
    .Q_t(n1859_t)
  );


  i1s3
  U4419
  (
    .DIN(n5110),
    .DIN_t(n5110_t),
    .Q(n1860),
    .Q_t(n1860_t)
  );


  i1s3
  U4420
  (
    .DIN(n5106),
    .DIN_t(n5106_t),
    .Q(n1861),
    .Q_t(n1861_t)
  );


  i1s3
  U4421
  (
    .DIN(n5102),
    .DIN_t(n5102_t),
    .Q(n1862),
    .Q_t(n1862_t)
  );


  i1s3
  U4422
  (
    .DIN(n5098),
    .DIN_t(n5098_t),
    .Q(n1863),
    .Q_t(n1863_t)
  );


  i1s3
  U4423
  (
    .DIN(n5094),
    .DIN_t(n5094_t),
    .Q(n1864),
    .Q_t(n1864_t)
  );


  i1s3
  U4424
  (
    .DIN(n5090),
    .DIN_t(n5090_t),
    .Q(n1865),
    .Q_t(n1865_t)
  );


  i1s3
  U4425
  (
    .DIN(n5086),
    .DIN_t(n5086_t),
    .Q(n1866),
    .Q_t(n1866_t)
  );


  i1s3
  U4426
  (
    .DIN(n5082),
    .DIN_t(n5082_t),
    .Q(n1867),
    .Q_t(n1867_t)
  );


  i1s3
  U4427
  (
    .DIN(n5078),
    .DIN_t(n5078_t),
    .Q(n1868),
    .Q_t(n1868_t)
  );


  i1s3
  U4428
  (
    .DIN(n5074),
    .DIN_t(n5074_t),
    .Q(n1869),
    .Q_t(n1869_t)
  );


  i1s3
  U4429
  (
    .DIN(n5070),
    .DIN_t(n5070_t),
    .Q(n1870),
    .Q_t(n1870_t)
  );


  i1s3
  U4430
  (
    .DIN(n5066),
    .DIN_t(n5066_t),
    .Q(n1871),
    .Q_t(n1871_t)
  );


  i1s3
  U4431
  (
    .DIN(n5062),
    .DIN_t(n5062_t),
    .Q(n1872),
    .Q_t(n1872_t)
  );


  i1s3
  U4432
  (
    .DIN(n5058),
    .DIN_t(n5058_t),
    .Q(n1873),
    .Q_t(n1873_t)
  );


  i1s3
  U4433
  (
    .DIN(n5054),
    .DIN_t(n5054_t),
    .Q(n1874),
    .Q_t(n1874_t)
  );


  i1s3
  U4434
  (
    .DIN(n5050),
    .DIN_t(n5050_t),
    .Q(n1875),
    .Q_t(n1875_t)
  );


  i1s3
  U4435
  (
    .DIN(n5046),
    .DIN_t(n5046_t),
    .Q(n1876),
    .Q_t(n1876_t)
  );


  i1s3
  U4436
  (
    .DIN(n5042),
    .DIN_t(n5042_t),
    .Q(n1877),
    .Q_t(n1877_t)
  );


  i1s3
  U4437
  (
    .DIN(n5038),
    .DIN_t(n5038_t),
    .Q(n1878),
    .Q_t(n1878_t)
  );


  i1s3
  U4438
  (
    .DIN(n5034),
    .DIN_t(n5034_t),
    .Q(n1879),
    .Q_t(n1879_t)
  );


  i1s3
  U4439
  (
    .DIN(n5030),
    .DIN_t(n5030_t),
    .Q(n1880),
    .Q_t(n1880_t)
  );


  i1s3
  U4440
  (
    .DIN(n5026),
    .DIN_t(n5026_t),
    .Q(n1881),
    .Q_t(n1881_t)
  );


  i1s3
  U4441
  (
    .DIN(n5022),
    .DIN_t(n5022_t),
    .Q(n1882),
    .Q_t(n1882_t)
  );


  i1s3
  U4442
  (
    .DIN(n5018),
    .DIN_t(n5018_t),
    .Q(n1883),
    .Q_t(n1883_t)
  );


  i1s3
  U4443
  (
    .DIN(n5014),
    .DIN_t(n5014_t),
    .Q(n1884),
    .Q_t(n1884_t)
  );


  i1s3
  U4444
  (
    .DIN(n5010),
    .DIN_t(n5010_t),
    .Q(n1885),
    .Q_t(n1885_t)
  );


  i1s3
  U4445
  (
    .DIN(n5006),
    .DIN_t(n5006_t),
    .Q(n1886),
    .Q_t(n1886_t)
  );


  i1s3
  U4446
  (
    .DIN(n5002),
    .DIN_t(n5002_t),
    .Q(n1887),
    .Q_t(n1887_t)
  );


  i1s3
  U4447
  (
    .DIN(n4998),
    .DIN_t(n4998_t),
    .Q(n1888),
    .Q_t(n1888_t)
  );


  i1s3
  U4448
  (
    .DIN(n5124),
    .DIN_t(n5124_t),
    .Q(n1889),
    .Q_t(n1889_t)
  );


  i1s3
  U4449
  (
    .DIN(n5125),
    .DIN_t(n5125_t),
    .Q(n1890),
    .Q_t(n1890_t)
  );


  i1s3
  U4450
  (
    .DIN(n5126),
    .DIN_t(n5126_t),
    .Q(n1891),
    .Q_t(n1891_t)
  );


  i1s3
  U4451
  (
    .DIN(n5127),
    .DIN_t(n5127_t),
    .Q(n1892),
    .Q_t(n1892_t)
  );


  i1s3
  U4452
  (
    .DIN(n5128),
    .DIN_t(n5128_t),
    .Q(n1893),
    .Q_t(n1893_t)
  );


  i1s3
  U4453
  (
    .DIN(n5129),
    .DIN_t(n5129_t),
    .Q(n1894),
    .Q_t(n1894_t)
  );


  i1s3
  U4454
  (
    .DIN(n5130),
    .DIN_t(n5130_t),
    .Q(n1895),
    .Q_t(n1895_t)
  );


  i1s3
  U4455
  (
    .DIN(n5131),
    .DIN_t(n5131_t),
    .Q(n1896),
    .Q_t(n1896_t)
  );


  i1s3
  U4456
  (
    .DIN(n5132),
    .DIN_t(n5132_t),
    .Q(n1897),
    .Q_t(n1897_t)
  );


  i1s3
  U4457
  (
    .DIN(n5133),
    .DIN_t(n5133_t),
    .Q(n1898),
    .Q_t(n1898_t)
  );


  i1s3
  U4458
  (
    .DIN(n5134),
    .DIN_t(n5134_t),
    .Q(n1899),
    .Q_t(n1899_t)
  );


  i1s3
  U4459
  (
    .DIN(n5135),
    .DIN_t(n5135_t),
    .Q(n1900),
    .Q_t(n1900_t)
  );


  i1s3
  U4460
  (
    .DIN(n5136),
    .DIN_t(n5136_t),
    .Q(n1901),
    .Q_t(n1901_t)
  );


  i1s3
  U4461
  (
    .DIN(n5137),
    .DIN_t(n5137_t),
    .Q(n1902),
    .Q_t(n1902_t)
  );


  i1s3
  U4462
  (
    .DIN(n5138),
    .DIN_t(n5138_t),
    .Q(n1903),
    .Q_t(n1903_t)
  );


  i1s3
  U4463
  (
    .DIN(n5139),
    .DIN_t(n5139_t),
    .Q(n1904),
    .Q_t(n1904_t)
  );


  i1s3
  U4464
  (
    .DIN(n5140),
    .DIN_t(n5140_t),
    .Q(n1905),
    .Q_t(n1905_t)
  );


  i1s3
  U4465
  (
    .DIN(n5141),
    .DIN_t(n5141_t),
    .Q(n1906),
    .Q_t(n1906_t)
  );


  i1s3
  U4466
  (
    .DIN(n5142),
    .DIN_t(n5142_t),
    .Q(n1907),
    .Q_t(n1907_t)
  );


  i1s3
  U4467
  (
    .DIN(n5143),
    .DIN_t(n5143_t),
    .Q(n1908),
    .Q_t(n1908_t)
  );


  i1s3
  U4468
  (
    .DIN(n5144),
    .DIN_t(n5144_t),
    .Q(n1909),
    .Q_t(n1909_t)
  );


  i1s3
  U4469
  (
    .DIN(n5145),
    .DIN_t(n5145_t),
    .Q(n1910),
    .Q_t(n1910_t)
  );


  i1s3
  U4470
  (
    .DIN(n5146),
    .DIN_t(n5146_t),
    .Q(n1911),
    .Q_t(n1911_t)
  );


  i1s3
  U4471
  (
    .DIN(n5147),
    .DIN_t(n5147_t),
    .Q(n1912),
    .Q_t(n1912_t)
  );


  i1s3
  U4472
  (
    .DIN(n5148),
    .DIN_t(n5148_t),
    .Q(n1913),
    .Q_t(n1913_t)
  );


  i1s3
  U4473
  (
    .DIN(n5149),
    .DIN_t(n5149_t),
    .Q(n1914),
    .Q_t(n1914_t)
  );


  i1s3
  U4474
  (
    .DIN(n5150),
    .DIN_t(n5150_t),
    .Q(n1915),
    .Q_t(n1915_t)
  );


  i1s3
  U4475
  (
    .DIN(n5151),
    .DIN_t(n5151_t),
    .Q(n1916),
    .Q_t(n1916_t)
  );


  i1s3
  U4476
  (
    .DIN(n5152),
    .DIN_t(n5152_t),
    .Q(n1917),
    .Q_t(n1917_t)
  );


  i1s3
  U4477
  (
    .DIN(n5153),
    .DIN_t(n5153_t),
    .Q(n1918),
    .Q_t(n1918_t)
  );


  i1s3
  U4478
  (
    .DIN(n5154),
    .DIN_t(n5154_t),
    .Q(n1919),
    .Q_t(n1919_t)
  );


  i1s3
  U4479
  (
    .DIN(n5123),
    .DIN_t(n5123_t),
    .Q(n1920),
    .Q_t(n1920_t)
  );


  i1s3
  U4480
  (
    .DIN(n5298),
    .DIN_t(n5298_t),
    .Q(n1921),
    .Q_t(n1921_t)
  );


  i1s3
  U4481
  (
    .DIN(n5293),
    .DIN_t(n5293_t),
    .Q(n1922),
    .Q_t(n1922_t)
  );


  i1s3
  U4482
  (
    .DIN(n5288),
    .DIN_t(n5288_t),
    .Q(n1923),
    .Q_t(n1923_t)
  );


  i1s3
  U4483
  (
    .DIN(n5283),
    .DIN_t(n5283_t),
    .Q(n1924),
    .Q_t(n1924_t)
  );


  i1s3
  U4484
  (
    .DIN(n5278),
    .DIN_t(n5278_t),
    .Q(n1925),
    .Q_t(n1925_t)
  );


  i1s3
  U4485
  (
    .DIN(n5273),
    .DIN_t(n5273_t),
    .Q(n1926),
    .Q_t(n1926_t)
  );


  i1s3
  U4486
  (
    .DIN(n5268),
    .DIN_t(n5268_t),
    .Q(n1927),
    .Q_t(n1927_t)
  );


  i1s3
  U4487
  (
    .DIN(n5263),
    .DIN_t(n5263_t),
    .Q(n1928),
    .Q_t(n1928_t)
  );


  i1s3
  U4488
  (
    .DIN(n5258),
    .DIN_t(n5258_t),
    .Q(n1929),
    .Q_t(n1929_t)
  );


  i1s3
  U4489
  (
    .DIN(n5253),
    .DIN_t(n5253_t),
    .Q(n1930),
    .Q_t(n1930_t)
  );


  i1s3
  U4490
  (
    .DIN(n5248),
    .DIN_t(n5248_t),
    .Q(n1931),
    .Q_t(n1931_t)
  );


  i1s3
  U4491
  (
    .DIN(n5243),
    .DIN_t(n5243_t),
    .Q(n1932),
    .Q_t(n1932_t)
  );


  i1s3
  U4492
  (
    .DIN(n5238),
    .DIN_t(n5238_t),
    .Q(n1933),
    .Q_t(n1933_t)
  );


  i1s3
  U4493
  (
    .DIN(n5233),
    .DIN_t(n5233_t),
    .Q(n1934),
    .Q_t(n1934_t)
  );


  i1s3
  U4494
  (
    .DIN(n5228),
    .DIN_t(n5228_t),
    .Q(n1935),
    .Q_t(n1935_t)
  );


  i1s3
  U4495
  (
    .DIN(n5223),
    .DIN_t(n5223_t),
    .Q(n1936),
    .Q_t(n1936_t)
  );


  i1s3
  U4496
  (
    .DIN(n5218),
    .DIN_t(n5218_t),
    .Q(n1937),
    .Q_t(n1937_t)
  );


  i1s3
  U4497
  (
    .DIN(n5214),
    .DIN_t(n5214_t),
    .Q(n1938),
    .Q_t(n1938_t)
  );


  i1s3
  U4498
  (
    .DIN(n5210),
    .DIN_t(n5210_t),
    .Q(n1939),
    .Q_t(n1939_t)
  );


  i1s3
  U4499
  (
    .DIN(n5206),
    .DIN_t(n5206_t),
    .Q(n1940),
    .Q_t(n1940_t)
  );


  i1s3
  U4500
  (
    .DIN(n5202),
    .DIN_t(n5202_t),
    .Q(n1941),
    .Q_t(n1941_t)
  );


  i1s3
  U4501
  (
    .DIN(n5198),
    .DIN_t(n5198_t),
    .Q(n1942),
    .Q_t(n1942_t)
  );


  i1s3
  U4502
  (
    .DIN(n5194),
    .DIN_t(n5194_t),
    .Q(n1943),
    .Q_t(n1943_t)
  );


  i1s3
  U4503
  (
    .DIN(n5190),
    .DIN_t(n5190_t),
    .Q(n1944),
    .Q_t(n1944_t)
  );


  i1s3
  U4504
  (
    .DIN(n5186),
    .DIN_t(n5186_t),
    .Q(n1945),
    .Q_t(n1945_t)
  );


  i1s3
  U4505
  (
    .DIN(n5182),
    .DIN_t(n5182_t),
    .Q(n1946),
    .Q_t(n1946_t)
  );


  i1s3
  U4506
  (
    .DIN(n5178),
    .DIN_t(n5178_t),
    .Q(n1947),
    .Q_t(n1947_t)
  );


  i1s3
  U4507
  (
    .DIN(n5174),
    .DIN_t(n5174_t),
    .Q(n1948),
    .Q_t(n1948_t)
  );


  i1s3
  U4508
  (
    .DIN(n5170),
    .DIN_t(n5170_t),
    .Q(n1949),
    .Q_t(n1949_t)
  );


  i1s3
  U4509
  (
    .DIN(n5166),
    .DIN_t(n5166_t),
    .Q(n1950),
    .Q_t(n1950_t)
  );


  i1s3
  U4510
  (
    .DIN(n5162),
    .DIN_t(n5162_t),
    .Q(n1951),
    .Q_t(n1951_t)
  );


  i1s3
  U4511
  (
    .DIN(n5158),
    .DIN_t(n5158_t),
    .Q(n1952),
    .Q_t(n1952_t)
  );


  i1s3
  U4512
  (
    .DIN(n5300),
    .DIN_t(n5300_t),
    .Q(n1953),
    .Q_t(n1953_t)
  );


  i1s3
  U4513
  (
    .DIN(n5301),
    .DIN_t(n5301_t),
    .Q(n1954),
    .Q_t(n1954_t)
  );


  i1s3
  U4514
  (
    .DIN(n5302),
    .DIN_t(n5302_t),
    .Q(n1955),
    .Q_t(n1955_t)
  );


  i1s3
  U4515
  (
    .DIN(n5303),
    .DIN_t(n5303_t),
    .Q(n1956),
    .Q_t(n1956_t)
  );


  i1s3
  U4516
  (
    .DIN(n5304),
    .DIN_t(n5304_t),
    .Q(n1957),
    .Q_t(n1957_t)
  );


  i1s3
  U4517
  (
    .DIN(n5305),
    .DIN_t(n5305_t),
    .Q(n1958),
    .Q_t(n1958_t)
  );


  i1s3
  U4518
  (
    .DIN(n5306),
    .DIN_t(n5306_t),
    .Q(n1959),
    .Q_t(n1959_t)
  );


  i1s3
  U4519
  (
    .DIN(n5307),
    .DIN_t(n5307_t),
    .Q(n1960),
    .Q_t(n1960_t)
  );


  i1s3
  U4520
  (
    .DIN(n5308),
    .DIN_t(n5308_t),
    .Q(n1961),
    .Q_t(n1961_t)
  );


  i1s3
  U4521
  (
    .DIN(n5309),
    .DIN_t(n5309_t),
    .Q(n1962),
    .Q_t(n1962_t)
  );


  i1s3
  U4522
  (
    .DIN(n5310),
    .DIN_t(n5310_t),
    .Q(n1963),
    .Q_t(n1963_t)
  );


  i1s3
  U4523
  (
    .DIN(n5311),
    .DIN_t(n5311_t),
    .Q(n1964),
    .Q_t(n1964_t)
  );


  i1s3
  U4524
  (
    .DIN(n5312),
    .DIN_t(n5312_t),
    .Q(n1965),
    .Q_t(n1965_t)
  );


  i1s3
  U4525
  (
    .DIN(n5313),
    .DIN_t(n5313_t),
    .Q(n1966),
    .Q_t(n1966_t)
  );


  i1s3
  U4526
  (
    .DIN(n5314),
    .DIN_t(n5314_t),
    .Q(n1967),
    .Q_t(n1967_t)
  );


  i1s3
  U4527
  (
    .DIN(n5315),
    .DIN_t(n5315_t),
    .Q(n1968),
    .Q_t(n1968_t)
  );


  i1s3
  U4528
  (
    .DIN(n5316),
    .DIN_t(n5316_t),
    .Q(n1969),
    .Q_t(n1969_t)
  );


  i1s3
  U4529
  (
    .DIN(n5317),
    .DIN_t(n5317_t),
    .Q(n1970),
    .Q_t(n1970_t)
  );


  i1s3
  U4530
  (
    .DIN(n5318),
    .DIN_t(n5318_t),
    .Q(n1971),
    .Q_t(n1971_t)
  );


  i1s3
  U4531
  (
    .DIN(n5319),
    .DIN_t(n5319_t),
    .Q(n1972),
    .Q_t(n1972_t)
  );


  i1s3
  U4532
  (
    .DIN(n5320),
    .DIN_t(n5320_t),
    .Q(n1973),
    .Q_t(n1973_t)
  );


  i1s3
  U4533
  (
    .DIN(n5321),
    .DIN_t(n5321_t),
    .Q(n1974),
    .Q_t(n1974_t)
  );


  i1s3
  U4534
  (
    .DIN(n5322),
    .DIN_t(n5322_t),
    .Q(n1975),
    .Q_t(n1975_t)
  );


  i1s3
  U4535
  (
    .DIN(n5323),
    .DIN_t(n5323_t),
    .Q(n1976),
    .Q_t(n1976_t)
  );


  i1s3
  U4536
  (
    .DIN(n5324),
    .DIN_t(n5324_t),
    .Q(n1977),
    .Q_t(n1977_t)
  );


  i1s3
  U4537
  (
    .DIN(n5325),
    .DIN_t(n5325_t),
    .Q(n1978),
    .Q_t(n1978_t)
  );


  i1s3
  U4538
  (
    .DIN(n5326),
    .DIN_t(n5326_t),
    .Q(n1979),
    .Q_t(n1979_t)
  );


  i1s3
  U4539
  (
    .DIN(n5327),
    .DIN_t(n5327_t),
    .Q(n1980),
    .Q_t(n1980_t)
  );


  i1s3
  U4540
  (
    .DIN(n5328),
    .DIN_t(n5328_t),
    .Q(n1981),
    .Q_t(n1981_t)
  );


  i1s3
  U4541
  (
    .DIN(n5329),
    .DIN_t(n5329_t),
    .Q(n1982),
    .Q_t(n1982_t)
  );


  i1s3
  U4542
  (
    .DIN(n5330),
    .DIN_t(n5330_t),
    .Q(n1983),
    .Q_t(n1983_t)
  );


  i1s3
  U4543
  (
    .DIN(n5299),
    .DIN_t(n5299_t),
    .Q(n1984),
    .Q_t(n1984_t)
  );


  i1s3
  U4544
  (
    .DIN(n5474),
    .DIN_t(n5474_t),
    .Q(n1985),
    .Q_t(n1985_t)
  );


  i1s3
  U4545
  (
    .DIN(n5469),
    .DIN_t(n5469_t),
    .Q(n1986),
    .Q_t(n1986_t)
  );


  i1s3
  U4546
  (
    .DIN(n5464),
    .DIN_t(n5464_t),
    .Q(n1987),
    .Q_t(n1987_t)
  );


  i1s3
  U4547
  (
    .DIN(n5459),
    .DIN_t(n5459_t),
    .Q(n1988),
    .Q_t(n1988_t)
  );


  i1s3
  U4548
  (
    .DIN(n5454),
    .DIN_t(n5454_t),
    .Q(n1989),
    .Q_t(n1989_t)
  );


  i1s3
  U4549
  (
    .DIN(n5449),
    .DIN_t(n5449_t),
    .Q(n1990),
    .Q_t(n1990_t)
  );


  i1s3
  U4550
  (
    .DIN(n5444),
    .DIN_t(n5444_t),
    .Q(n1991),
    .Q_t(n1991_t)
  );


  i1s3
  U4551
  (
    .DIN(n5439),
    .DIN_t(n5439_t),
    .Q(n1992),
    .Q_t(n1992_t)
  );


  i1s3
  U4552
  (
    .DIN(n5434),
    .DIN_t(n5434_t),
    .Q(n1993),
    .Q_t(n1993_t)
  );


  i1s3
  U4553
  (
    .DIN(n5429),
    .DIN_t(n5429_t),
    .Q(n1994),
    .Q_t(n1994_t)
  );


  i1s3
  U4554
  (
    .DIN(n5424),
    .DIN_t(n5424_t),
    .Q(n1995),
    .Q_t(n1995_t)
  );


  i1s3
  U4555
  (
    .DIN(n5419),
    .DIN_t(n5419_t),
    .Q(n1996),
    .Q_t(n1996_t)
  );


  i1s3
  U4556
  (
    .DIN(n5414),
    .DIN_t(n5414_t),
    .Q(n1997),
    .Q_t(n1997_t)
  );


  i1s3
  U4557
  (
    .DIN(n5409),
    .DIN_t(n5409_t),
    .Q(n1998),
    .Q_t(n1998_t)
  );


  i1s3
  U4558
  (
    .DIN(n5404),
    .DIN_t(n5404_t),
    .Q(n1999),
    .Q_t(n1999_t)
  );


  i1s3
  U4559
  (
    .DIN(n5399),
    .DIN_t(n5399_t),
    .Q(n2000),
    .Q_t(n2000_t)
  );


  i1s3
  U4560
  (
    .DIN(n5394),
    .DIN_t(n5394_t),
    .Q(n2001),
    .Q_t(n2001_t)
  );


  i1s3
  U4561
  (
    .DIN(n5390),
    .DIN_t(n5390_t),
    .Q(n2002),
    .Q_t(n2002_t)
  );


  i1s3
  U4562
  (
    .DIN(n5386),
    .DIN_t(n5386_t),
    .Q(n2003),
    .Q_t(n2003_t)
  );


  i1s3
  U4563
  (
    .DIN(n5382),
    .DIN_t(n5382_t),
    .Q(n2004),
    .Q_t(n2004_t)
  );


  i1s3
  U4564
  (
    .DIN(n5378),
    .DIN_t(n5378_t),
    .Q(n2005),
    .Q_t(n2005_t)
  );


  i1s3
  U4565
  (
    .DIN(n5374),
    .DIN_t(n5374_t),
    .Q(n2006),
    .Q_t(n2006_t)
  );


  i1s3
  U4566
  (
    .DIN(n5370),
    .DIN_t(n5370_t),
    .Q(n2007),
    .Q_t(n2007_t)
  );


  i1s3
  U4567
  (
    .DIN(n5366),
    .DIN_t(n5366_t),
    .Q(n2008),
    .Q_t(n2008_t)
  );


  i1s3
  U4568
  (
    .DIN(n5362),
    .DIN_t(n5362_t),
    .Q(n2009),
    .Q_t(n2009_t)
  );


  i1s3
  U4569
  (
    .DIN(n5358),
    .DIN_t(n5358_t),
    .Q(n2010),
    .Q_t(n2010_t)
  );


  i1s3
  U4570
  (
    .DIN(n5354),
    .DIN_t(n5354_t),
    .Q(n2011),
    .Q_t(n2011_t)
  );


  i1s3
  U4571
  (
    .DIN(n5350),
    .DIN_t(n5350_t),
    .Q(n2012),
    .Q_t(n2012_t)
  );


  i1s3
  U4572
  (
    .DIN(n5346),
    .DIN_t(n5346_t),
    .Q(n2013),
    .Q_t(n2013_t)
  );


  i1s3
  U4573
  (
    .DIN(n5342),
    .DIN_t(n5342_t),
    .Q(n2014),
    .Q_t(n2014_t)
  );


  i1s3
  U4574
  (
    .DIN(n5338),
    .DIN_t(n5338_t),
    .Q(n2015),
    .Q_t(n2015_t)
  );


  i1s3
  U4575
  (
    .DIN(n5334),
    .DIN_t(n5334_t),
    .Q(n2016),
    .Q_t(n2016_t)
  );


  i1s3
  U4576
  (
    .DIN(n5476),
    .DIN_t(n5476_t),
    .Q(n2017),
    .Q_t(n2017_t)
  );


  i1s3
  U4577
  (
    .DIN(n5477),
    .DIN_t(n5477_t),
    .Q(n2018),
    .Q_t(n2018_t)
  );


  i1s3
  U4578
  (
    .DIN(n5478),
    .DIN_t(n5478_t),
    .Q(n2019),
    .Q_t(n2019_t)
  );


  i1s3
  U4579
  (
    .DIN(n5479),
    .DIN_t(n5479_t),
    .Q(n2020),
    .Q_t(n2020_t)
  );


  i1s3
  U4580
  (
    .DIN(n5480),
    .DIN_t(n5480_t),
    .Q(n2021),
    .Q_t(n2021_t)
  );


  i1s3
  U4581
  (
    .DIN(n5481),
    .DIN_t(n5481_t),
    .Q(n2022),
    .Q_t(n2022_t)
  );


  i1s3
  U4582
  (
    .DIN(n5482),
    .DIN_t(n5482_t),
    .Q(n2023),
    .Q_t(n2023_t)
  );


  i1s3
  U4583
  (
    .DIN(n5483),
    .DIN_t(n5483_t),
    .Q(n2024),
    .Q_t(n2024_t)
  );


  i1s3
  U4584
  (
    .DIN(n5484),
    .DIN_t(n5484_t),
    .Q(n2025),
    .Q_t(n2025_t)
  );


  i1s3
  U4585
  (
    .DIN(n5485),
    .DIN_t(n5485_t),
    .Q(n2026),
    .Q_t(n2026_t)
  );


  i1s3
  U4586
  (
    .DIN(n5486),
    .DIN_t(n5486_t),
    .Q(n2027),
    .Q_t(n2027_t)
  );


  i1s3
  U4587
  (
    .DIN(n5487),
    .DIN_t(n5487_t),
    .Q(n2028),
    .Q_t(n2028_t)
  );


  i1s3
  U4588
  (
    .DIN(n5488),
    .DIN_t(n5488_t),
    .Q(n2029),
    .Q_t(n2029_t)
  );


  i1s3
  U4589
  (
    .DIN(n5489),
    .DIN_t(n5489_t),
    .Q(n2030),
    .Q_t(n2030_t)
  );


  i1s3
  U4590
  (
    .DIN(n5490),
    .DIN_t(n5490_t),
    .Q(n2031),
    .Q_t(n2031_t)
  );


  i1s3
  U4591
  (
    .DIN(n5491),
    .DIN_t(n5491_t),
    .Q(n2032),
    .Q_t(n2032_t)
  );


  i1s3
  U4592
  (
    .DIN(n5492),
    .DIN_t(n5492_t),
    .Q(n2033),
    .Q_t(n2033_t)
  );


  i1s3
  U4593
  (
    .DIN(n5493),
    .DIN_t(n5493_t),
    .Q(n2034),
    .Q_t(n2034_t)
  );


  i1s3
  U4594
  (
    .DIN(n5494),
    .DIN_t(n5494_t),
    .Q(n2035),
    .Q_t(n2035_t)
  );


  i1s3
  U4595
  (
    .DIN(n5495),
    .DIN_t(n5495_t),
    .Q(n2036),
    .Q_t(n2036_t)
  );


  i1s3
  U4596
  (
    .DIN(n5496),
    .DIN_t(n5496_t),
    .Q(n2037),
    .Q_t(n2037_t)
  );


  i1s3
  U4597
  (
    .DIN(n5497),
    .DIN_t(n5497_t),
    .Q(n2038),
    .Q_t(n2038_t)
  );


  i1s3
  U4598
  (
    .DIN(n5498),
    .DIN_t(n5498_t),
    .Q(n2039),
    .Q_t(n2039_t)
  );


  i1s3
  U4599
  (
    .DIN(n5499),
    .DIN_t(n5499_t),
    .Q(n2040),
    .Q_t(n2040_t)
  );


  i1s3
  U4600
  (
    .DIN(n5500),
    .DIN_t(n5500_t),
    .Q(n2041),
    .Q_t(n2041_t)
  );


  i1s3
  U4601
  (
    .DIN(n5501),
    .DIN_t(n5501_t),
    .Q(n2042),
    .Q_t(n2042_t)
  );


  i1s3
  U4602
  (
    .DIN(n5502),
    .DIN_t(n5502_t),
    .Q(n2043),
    .Q_t(n2043_t)
  );


  i1s3
  U4603
  (
    .DIN(n5503),
    .DIN_t(n5503_t),
    .Q(n2044),
    .Q_t(n2044_t)
  );


  i1s3
  U4604
  (
    .DIN(n5504),
    .DIN_t(n5504_t),
    .Q(n2045),
    .Q_t(n2045_t)
  );


  i1s3
  U4605
  (
    .DIN(n5505),
    .DIN_t(n5505_t),
    .Q(n2046),
    .Q_t(n2046_t)
  );


  i1s3
  U4606
  (
    .DIN(n5506),
    .DIN_t(n5506_t),
    .Q(n2047),
    .Q_t(n2047_t)
  );


  i1s3
  U4607
  (
    .DIN(n5475),
    .DIN_t(n5475_t),
    .Q(n2048),
    .Q_t(n2048_t)
  );


  i1s3
  U4608
  (
    .DIN(n5650),
    .DIN_t(n5650_t),
    .Q(n2049),
    .Q_t(n2049_t)
  );


  i1s3
  U4609
  (
    .DIN(n5645),
    .DIN_t(n5645_t),
    .Q(n2050),
    .Q_t(n2050_t)
  );


  i1s3
  U4610
  (
    .DIN(n5640),
    .DIN_t(n5640_t),
    .Q(n2051),
    .Q_t(n2051_t)
  );


  i1s3
  U4611
  (
    .DIN(n5635),
    .DIN_t(n5635_t),
    .Q(n2052),
    .Q_t(n2052_t)
  );


  i1s3
  U4612
  (
    .DIN(n5630),
    .DIN_t(n5630_t),
    .Q(n2053),
    .Q_t(n2053_t)
  );


  i1s3
  U4613
  (
    .DIN(n5625),
    .DIN_t(n5625_t),
    .Q(n2054),
    .Q_t(n2054_t)
  );


  i1s3
  U4614
  (
    .DIN(n5620),
    .DIN_t(n5620_t),
    .Q(n2055),
    .Q_t(n2055_t)
  );


  i1s3
  U4615
  (
    .DIN(n5615),
    .DIN_t(n5615_t),
    .Q(n2056),
    .Q_t(n2056_t)
  );


  i1s3
  U4616
  (
    .DIN(n5610),
    .DIN_t(n5610_t),
    .Q(n2057),
    .Q_t(n2057_t)
  );


  i1s3
  U4617
  (
    .DIN(n5605),
    .DIN_t(n5605_t),
    .Q(n2058),
    .Q_t(n2058_t)
  );


  i1s3
  U4618
  (
    .DIN(n5600),
    .DIN_t(n5600_t),
    .Q(n2059),
    .Q_t(n2059_t)
  );


  i1s3
  U4619
  (
    .DIN(n5595),
    .DIN_t(n5595_t),
    .Q(n2060),
    .Q_t(n2060_t)
  );


  i1s3
  U4620
  (
    .DIN(n5590),
    .DIN_t(n5590_t),
    .Q(n2061),
    .Q_t(n2061_t)
  );


  i1s3
  U4621
  (
    .DIN(n5585),
    .DIN_t(n5585_t),
    .Q(n2062),
    .Q_t(n2062_t)
  );


  i1s3
  U4622
  (
    .DIN(n5580),
    .DIN_t(n5580_t),
    .Q(n2063),
    .Q_t(n2063_t)
  );


  i1s3
  U4623
  (
    .DIN(n5575),
    .DIN_t(n5575_t),
    .Q(n2064),
    .Q_t(n2064_t)
  );


  i1s3
  U4624
  (
    .DIN(n5570),
    .DIN_t(n5570_t),
    .Q(n2065),
    .Q_t(n2065_t)
  );


  i1s3
  U4625
  (
    .DIN(n5566),
    .DIN_t(n5566_t),
    .Q(n2066),
    .Q_t(n2066_t)
  );


  i1s3
  U4626
  (
    .DIN(n5562),
    .DIN_t(n5562_t),
    .Q(n2067),
    .Q_t(n2067_t)
  );


  i1s3
  U4627
  (
    .DIN(n5558),
    .DIN_t(n5558_t),
    .Q(n2068),
    .Q_t(n2068_t)
  );


  i1s3
  U4628
  (
    .DIN(n5554),
    .DIN_t(n5554_t),
    .Q(n2069),
    .Q_t(n2069_t)
  );


  i1s3
  U4629
  (
    .DIN(n5550),
    .DIN_t(n5550_t),
    .Q(n2070),
    .Q_t(n2070_t)
  );


  i1s3
  U4630
  (
    .DIN(n5546),
    .DIN_t(n5546_t),
    .Q(n2071),
    .Q_t(n2071_t)
  );


  i1s3
  U4631
  (
    .DIN(n5542),
    .DIN_t(n5542_t),
    .Q(n2072),
    .Q_t(n2072_t)
  );


  i1s3
  U4632
  (
    .DIN(n5538),
    .DIN_t(n5538_t),
    .Q(n2073),
    .Q_t(n2073_t)
  );


  i1s3
  U4633
  (
    .DIN(n5534),
    .DIN_t(n5534_t),
    .Q(n2074),
    .Q_t(n2074_t)
  );


  i1s3
  U4634
  (
    .DIN(n5530),
    .DIN_t(n5530_t),
    .Q(n2075),
    .Q_t(n2075_t)
  );


  i1s3
  U4635
  (
    .DIN(n5526),
    .DIN_t(n5526_t),
    .Q(n2076),
    .Q_t(n2076_t)
  );


  i1s3
  U4636
  (
    .DIN(n5522),
    .DIN_t(n5522_t),
    .Q(n2077),
    .Q_t(n2077_t)
  );


  i1s3
  U4637
  (
    .DIN(n5518),
    .DIN_t(n5518_t),
    .Q(n2078),
    .Q_t(n2078_t)
  );


  i1s3
  U4638
  (
    .DIN(n5514),
    .DIN_t(n5514_t),
    .Q(n2079),
    .Q_t(n2079_t)
  );


  i1s3
  U4639
  (
    .DIN(n5510),
    .DIN_t(n5510_t),
    .Q(n2080),
    .Q_t(n2080_t)
  );


  i1s3
  U4640
  (
    .DIN(n5652),
    .DIN_t(n5652_t),
    .Q(n2081),
    .Q_t(n2081_t)
  );


  i1s3
  U4641
  (
    .DIN(n5653),
    .DIN_t(n5653_t),
    .Q(n2082),
    .Q_t(n2082_t)
  );


  i1s3
  U4642
  (
    .DIN(n5654),
    .DIN_t(n5654_t),
    .Q(n2083),
    .Q_t(n2083_t)
  );


  i1s3
  U4643
  (
    .DIN(n5655),
    .DIN_t(n5655_t),
    .Q(n2084),
    .Q_t(n2084_t)
  );


  i1s3
  U4644
  (
    .DIN(n5656),
    .DIN_t(n5656_t),
    .Q(n2085),
    .Q_t(n2085_t)
  );


  i1s3
  U4645
  (
    .DIN(n5657),
    .DIN_t(n5657_t),
    .Q(n2086),
    .Q_t(n2086_t)
  );


  i1s3
  U4646
  (
    .DIN(n5658),
    .DIN_t(n5658_t),
    .Q(n2087),
    .Q_t(n2087_t)
  );


  i1s3
  U4647
  (
    .DIN(n5659),
    .DIN_t(n5659_t),
    .Q(n2088),
    .Q_t(n2088_t)
  );


  i1s3
  U4648
  (
    .DIN(n5660),
    .DIN_t(n5660_t),
    .Q(n2089),
    .Q_t(n2089_t)
  );


  i1s3
  U4649
  (
    .DIN(n5661),
    .DIN_t(n5661_t),
    .Q(n2090),
    .Q_t(n2090_t)
  );


  i1s3
  U4650
  (
    .DIN(n5662),
    .DIN_t(n5662_t),
    .Q(n2091),
    .Q_t(n2091_t)
  );


  i1s3
  U4651
  (
    .DIN(n5663),
    .DIN_t(n5663_t),
    .Q(n2092),
    .Q_t(n2092_t)
  );


  i1s3
  U4652
  (
    .DIN(n5664),
    .DIN_t(n5664_t),
    .Q(n2093),
    .Q_t(n2093_t)
  );


  i1s3
  U4653
  (
    .DIN(n5665),
    .DIN_t(n5665_t),
    .Q(n2094),
    .Q_t(n2094_t)
  );


  i1s3
  U4654
  (
    .DIN(n5666),
    .DIN_t(n5666_t),
    .Q(n2095),
    .Q_t(n2095_t)
  );


  i1s3
  U4655
  (
    .DIN(n5667),
    .DIN_t(n5667_t),
    .Q(n2096),
    .Q_t(n2096_t)
  );


  i1s3
  U4656
  (
    .DIN(n5668),
    .DIN_t(n5668_t),
    .Q(n2097),
    .Q_t(n2097_t)
  );


  i1s3
  U4657
  (
    .DIN(n5669),
    .DIN_t(n5669_t),
    .Q(n2098),
    .Q_t(n2098_t)
  );


  i1s3
  U4658
  (
    .DIN(n5670),
    .DIN_t(n5670_t),
    .Q(n2099),
    .Q_t(n2099_t)
  );


  i1s3
  U4659
  (
    .DIN(n5671),
    .DIN_t(n5671_t),
    .Q(n2100),
    .Q_t(n2100_t)
  );


  i1s3
  U4660
  (
    .DIN(n5672),
    .DIN_t(n5672_t),
    .Q(n2101),
    .Q_t(n2101_t)
  );


  i1s3
  U4661
  (
    .DIN(n5673),
    .DIN_t(n5673_t),
    .Q(n2102),
    .Q_t(n2102_t)
  );


  i1s3
  U4662
  (
    .DIN(n5674),
    .DIN_t(n5674_t),
    .Q(n2103),
    .Q_t(n2103_t)
  );


  i1s3
  U4663
  (
    .DIN(n5675),
    .DIN_t(n5675_t),
    .Q(n2104),
    .Q_t(n2104_t)
  );


  i1s3
  U4664
  (
    .DIN(n5676),
    .DIN_t(n5676_t),
    .Q(n2105),
    .Q_t(n2105_t)
  );


  i1s3
  U4665
  (
    .DIN(n5677),
    .DIN_t(n5677_t),
    .Q(n2106),
    .Q_t(n2106_t)
  );


  i1s3
  U4666
  (
    .DIN(n5678),
    .DIN_t(n5678_t),
    .Q(n2107),
    .Q_t(n2107_t)
  );


  i1s3
  U4667
  (
    .DIN(n5679),
    .DIN_t(n5679_t),
    .Q(n2108),
    .Q_t(n2108_t)
  );


  i1s3
  U4668
  (
    .DIN(n5680),
    .DIN_t(n5680_t),
    .Q(n2109),
    .Q_t(n2109_t)
  );


  i1s3
  U4669
  (
    .DIN(n5681),
    .DIN_t(n5681_t),
    .Q(n2110),
    .Q_t(n2110_t)
  );


  i1s3
  U4670
  (
    .DIN(n5682),
    .DIN_t(n5682_t),
    .Q(n2111),
    .Q_t(n2111_t)
  );


  i1s3
  U4671
  (
    .DIN(n5651),
    .DIN_t(n5651_t),
    .Q(n2112),
    .Q_t(n2112_t)
  );


  i1s3
  U4672
  (
    .DIN(n5826),
    .DIN_t(n5826_t),
    .Q(n2113),
    .Q_t(n2113_t)
  );


  i1s3
  U4673
  (
    .DIN(n5821),
    .DIN_t(n5821_t),
    .Q(n2114),
    .Q_t(n2114_t)
  );


  i1s3
  U4674
  (
    .DIN(n5816),
    .DIN_t(n5816_t),
    .Q(n2115),
    .Q_t(n2115_t)
  );


  i1s3
  U4675
  (
    .DIN(n5811),
    .DIN_t(n5811_t),
    .Q(n2116),
    .Q_t(n2116_t)
  );


  i1s3
  U4676
  (
    .DIN(n5806),
    .DIN_t(n5806_t),
    .Q(n2117),
    .Q_t(n2117_t)
  );


  i1s3
  U4677
  (
    .DIN(n5801),
    .DIN_t(n5801_t),
    .Q(n2118),
    .Q_t(n2118_t)
  );


  i1s3
  U4678
  (
    .DIN(n5796),
    .DIN_t(n5796_t),
    .Q(n2119),
    .Q_t(n2119_t)
  );


  i1s3
  U4679
  (
    .DIN(n5791),
    .DIN_t(n5791_t),
    .Q(n2120),
    .Q_t(n2120_t)
  );


  i1s3
  U4680
  (
    .DIN(n5786),
    .DIN_t(n5786_t),
    .Q(n2121),
    .Q_t(n2121_t)
  );


  i1s3
  U4681
  (
    .DIN(n5781),
    .DIN_t(n5781_t),
    .Q(n2122),
    .Q_t(n2122_t)
  );


  i1s3
  U4682
  (
    .DIN(n5776),
    .DIN_t(n5776_t),
    .Q(n2123),
    .Q_t(n2123_t)
  );


  i1s3
  U4683
  (
    .DIN(n5771),
    .DIN_t(n5771_t),
    .Q(n2124),
    .Q_t(n2124_t)
  );


  i1s3
  U4684
  (
    .DIN(n5766),
    .DIN_t(n5766_t),
    .Q(n2125),
    .Q_t(n2125_t)
  );


  i1s3
  U4685
  (
    .DIN(n5761),
    .DIN_t(n5761_t),
    .Q(n2126),
    .Q_t(n2126_t)
  );


  i1s3
  U4686
  (
    .DIN(n5756),
    .DIN_t(n5756_t),
    .Q(n2127),
    .Q_t(n2127_t)
  );


  i1s3
  U4687
  (
    .DIN(n5751),
    .DIN_t(n5751_t),
    .Q(n2128),
    .Q_t(n2128_t)
  );


  i1s3
  U4688
  (
    .DIN(n5746),
    .DIN_t(n5746_t),
    .Q(n2129),
    .Q_t(n2129_t)
  );


  i1s3
  U4689
  (
    .DIN(n5742),
    .DIN_t(n5742_t),
    .Q(n2130),
    .Q_t(n2130_t)
  );


  i1s3
  U4690
  (
    .DIN(n5738),
    .DIN_t(n5738_t),
    .Q(n2131),
    .Q_t(n2131_t)
  );


  i1s3
  U4691
  (
    .DIN(n5734),
    .DIN_t(n5734_t),
    .Q(n2132),
    .Q_t(n2132_t)
  );


  i1s3
  U4692
  (
    .DIN(n5730),
    .DIN_t(n5730_t),
    .Q(n2133),
    .Q_t(n2133_t)
  );


  i1s3
  U4693
  (
    .DIN(n5726),
    .DIN_t(n5726_t),
    .Q(n2134),
    .Q_t(n2134_t)
  );


  i1s3
  U4694
  (
    .DIN(n5722),
    .DIN_t(n5722_t),
    .Q(n2135),
    .Q_t(n2135_t)
  );


  i1s3
  U4695
  (
    .DIN(n5718),
    .DIN_t(n5718_t),
    .Q(n2136),
    .Q_t(n2136_t)
  );


  i1s3
  U4696
  (
    .DIN(n5714),
    .DIN_t(n5714_t),
    .Q(n2137),
    .Q_t(n2137_t)
  );


  i1s3
  U4697
  (
    .DIN(n5710),
    .DIN_t(n5710_t),
    .Q(n2138),
    .Q_t(n2138_t)
  );


  i1s3
  U4698
  (
    .DIN(n5706),
    .DIN_t(n5706_t),
    .Q(n2139),
    .Q_t(n2139_t)
  );


  i1s3
  U4699
  (
    .DIN(n5702),
    .DIN_t(n5702_t),
    .Q(n2140),
    .Q_t(n2140_t)
  );


  i1s3
  U4700
  (
    .DIN(n5698),
    .DIN_t(n5698_t),
    .Q(n2141),
    .Q_t(n2141_t)
  );


  i1s3
  U4701
  (
    .DIN(n5694),
    .DIN_t(n5694_t),
    .Q(n2142),
    .Q_t(n2142_t)
  );


  i1s3
  U4702
  (
    .DIN(n5690),
    .DIN_t(n5690_t),
    .Q(n2143),
    .Q_t(n2143_t)
  );


  i1s3
  U4703
  (
    .DIN(n5686),
    .DIN_t(n5686_t),
    .Q(n2144),
    .Q_t(n2144_t)
  );


  i1s3
  U4704
  (
    .DIN(n5828),
    .DIN_t(n5828_t),
    .Q(n2145),
    .Q_t(n2145_t)
  );


  i1s3
  U4705
  (
    .DIN(n5829),
    .DIN_t(n5829_t),
    .Q(n2146),
    .Q_t(n2146_t)
  );


  i1s3
  U4706
  (
    .DIN(n5830),
    .DIN_t(n5830_t),
    .Q(n2147),
    .Q_t(n2147_t)
  );


  i1s3
  U4707
  (
    .DIN(n5831),
    .DIN_t(n5831_t),
    .Q(n2148),
    .Q_t(n2148_t)
  );


  i1s3
  U4708
  (
    .DIN(n5832),
    .DIN_t(n5832_t),
    .Q(n2149),
    .Q_t(n2149_t)
  );


  i1s3
  U4709
  (
    .DIN(n5833),
    .DIN_t(n5833_t),
    .Q(n2150),
    .Q_t(n2150_t)
  );


  i1s3
  U4710
  (
    .DIN(n5834),
    .DIN_t(n5834_t),
    .Q(n2151),
    .Q_t(n2151_t)
  );


  i1s3
  U4711
  (
    .DIN(n5835),
    .DIN_t(n5835_t),
    .Q(n2152),
    .Q_t(n2152_t)
  );


  i1s3
  U4712
  (
    .DIN(n5836),
    .DIN_t(n5836_t),
    .Q(n2153),
    .Q_t(n2153_t)
  );


  i1s3
  U4713
  (
    .DIN(n5837),
    .DIN_t(n5837_t),
    .Q(n2154),
    .Q_t(n2154_t)
  );


  i1s3
  U4714
  (
    .DIN(n5838),
    .DIN_t(n5838_t),
    .Q(n2155),
    .Q_t(n2155_t)
  );


  i1s3
  U4715
  (
    .DIN(n5839),
    .DIN_t(n5839_t),
    .Q(n2156),
    .Q_t(n2156_t)
  );


  i1s3
  U4716
  (
    .DIN(n5840),
    .DIN_t(n5840_t),
    .Q(n2157),
    .Q_t(n2157_t)
  );


  i1s3
  U4717
  (
    .DIN(n5841),
    .DIN_t(n5841_t),
    .Q(n2158),
    .Q_t(n2158_t)
  );


  i1s3
  U4718
  (
    .DIN(n5842),
    .DIN_t(n5842_t),
    .Q(n2159),
    .Q_t(n2159_t)
  );


  i1s3
  U4719
  (
    .DIN(n5843),
    .DIN_t(n5843_t),
    .Q(n2160),
    .Q_t(n2160_t)
  );


  i1s3
  U4720
  (
    .DIN(n5844),
    .DIN_t(n5844_t),
    .Q(n2161),
    .Q_t(n2161_t)
  );


  i1s3
  U4721
  (
    .DIN(n5845),
    .DIN_t(n5845_t),
    .Q(n2162),
    .Q_t(n2162_t)
  );


  i1s3
  U4722
  (
    .DIN(n5846),
    .DIN_t(n5846_t),
    .Q(n2163),
    .Q_t(n2163_t)
  );


  i1s3
  U4723
  (
    .DIN(n5847),
    .DIN_t(n5847_t),
    .Q(n2164),
    .Q_t(n2164_t)
  );


  i1s3
  U4724
  (
    .DIN(n5848),
    .DIN_t(n5848_t),
    .Q(n2165),
    .Q_t(n2165_t)
  );


  i1s3
  U4725
  (
    .DIN(n5849),
    .DIN_t(n5849_t),
    .Q(n2166),
    .Q_t(n2166_t)
  );


  i1s3
  U4726
  (
    .DIN(n5850),
    .DIN_t(n5850_t),
    .Q(n2167),
    .Q_t(n2167_t)
  );


  i1s3
  U4727
  (
    .DIN(n5851),
    .DIN_t(n5851_t),
    .Q(n2168),
    .Q_t(n2168_t)
  );


  i1s3
  U4728
  (
    .DIN(n5852),
    .DIN_t(n5852_t),
    .Q(n2169),
    .Q_t(n2169_t)
  );


  i1s3
  U4729
  (
    .DIN(n5853),
    .DIN_t(n5853_t),
    .Q(n2170),
    .Q_t(n2170_t)
  );


  i1s3
  U4730
  (
    .DIN(n5854),
    .DIN_t(n5854_t),
    .Q(n2171),
    .Q_t(n2171_t)
  );


  i1s3
  U4731
  (
    .DIN(n5855),
    .DIN_t(n5855_t),
    .Q(n2172),
    .Q_t(n2172_t)
  );


  i1s3
  U4732
  (
    .DIN(n5856),
    .DIN_t(n5856_t),
    .Q(n2173),
    .Q_t(n2173_t)
  );


  i1s3
  U4733
  (
    .DIN(n5857),
    .DIN_t(n5857_t),
    .Q(n2174),
    .Q_t(n2174_t)
  );


  i1s3
  U4734
  (
    .DIN(n5858),
    .DIN_t(n5858_t),
    .Q(n2175),
    .Q_t(n2175_t)
  );


  i1s3
  U4735
  (
    .DIN(n5827),
    .DIN_t(n5827_t),
    .Q(n2176),
    .Q_t(n2176_t)
  );


  i1s3
  U4736
  (
    .DIN(n6114),
    .DIN_t(n6114_t),
    .Q(n2177),
    .Q_t(n2177_t)
  );


  i1s3
  U4737
  (
    .DIN(n6105),
    .DIN_t(n6105_t),
    .Q(n2178),
    .Q_t(n2178_t)
  );


  i1s3
  U4738
  (
    .DIN(n6096),
    .DIN_t(n6096_t),
    .Q(n2179),
    .Q_t(n2179_t)
  );


  i1s3
  U4739
  (
    .DIN(n6087),
    .DIN_t(n6087_t),
    .Q(n2180),
    .Q_t(n2180_t)
  );


  i1s3
  U4740
  (
    .DIN(n6078),
    .DIN_t(n6078_t),
    .Q(n2181),
    .Q_t(n2181_t)
  );


  i1s3
  U4741
  (
    .DIN(n6069),
    .DIN_t(n6069_t),
    .Q(n2182),
    .Q_t(n2182_t)
  );


  i1s3
  U4742
  (
    .DIN(n6060),
    .DIN_t(n6060_t),
    .Q(n2183),
    .Q_t(n2183_t)
  );


  i1s3
  U4743
  (
    .DIN(n6051),
    .DIN_t(n6051_t),
    .Q(n2184),
    .Q_t(n2184_t)
  );


  i1s3
  U4744
  (
    .DIN(n6042),
    .DIN_t(n6042_t),
    .Q(n2185),
    .Q_t(n2185_t)
  );


  i1s3
  U4745
  (
    .DIN(n6033),
    .DIN_t(n6033_t),
    .Q(n2186),
    .Q_t(n2186_t)
  );


  i1s3
  U4746
  (
    .DIN(n6024),
    .DIN_t(n6024_t),
    .Q(n2187),
    .Q_t(n2187_t)
  );


  i1s3
  U4747
  (
    .DIN(n6015),
    .DIN_t(n6015_t),
    .Q(n2188),
    .Q_t(n2188_t)
  );


  i1s3
  U4748
  (
    .DIN(n6006),
    .DIN_t(n6006_t),
    .Q(n2189),
    .Q_t(n2189_t)
  );


  i1s3
  U4749
  (
    .DIN(n5997),
    .DIN_t(n5997_t),
    .Q(n2190),
    .Q_t(n2190_t)
  );


  i1s3
  U4750
  (
    .DIN(n5988),
    .DIN_t(n5988_t),
    .Q(n2191),
    .Q_t(n2191_t)
  );


  i1s3
  U4751
  (
    .DIN(n5979),
    .DIN_t(n5979_t),
    .Q(n2192),
    .Q_t(n2192_t)
  );


  i1s3
  U4752
  (
    .DIN(n5970),
    .DIN_t(n5970_t),
    .Q(n2193),
    .Q_t(n2193_t)
  );


  i1s3
  U4753
  (
    .DIN(n5963),
    .DIN_t(n5963_t),
    .Q(n2194),
    .Q_t(n2194_t)
  );


  i1s3
  U4754
  (
    .DIN(n5956),
    .DIN_t(n5956_t),
    .Q(n2195),
    .Q_t(n2195_t)
  );


  i1s3
  U4755
  (
    .DIN(n5949),
    .DIN_t(n5949_t),
    .Q(n2196),
    .Q_t(n2196_t)
  );


  i1s3
  U4756
  (
    .DIN(n5942),
    .DIN_t(n5942_t),
    .Q(n2197),
    .Q_t(n2197_t)
  );


  i1s3
  U4757
  (
    .DIN(n5935),
    .DIN_t(n5935_t),
    .Q(n2198),
    .Q_t(n2198_t)
  );


  i1s3
  U4758
  (
    .DIN(n5928),
    .DIN_t(n5928_t),
    .Q(n2199),
    .Q_t(n2199_t)
  );


  i1s3
  U4759
  (
    .DIN(n5921),
    .DIN_t(n5921_t),
    .Q(n2200),
    .Q_t(n2200_t)
  );


  i1s3
  U4760
  (
    .DIN(n5914),
    .DIN_t(n5914_t),
    .Q(n2201),
    .Q_t(n2201_t)
  );


  i1s3
  U4761
  (
    .DIN(n5907),
    .DIN_t(n5907_t),
    .Q(n2202),
    .Q_t(n2202_t)
  );


  i1s3
  U4762
  (
    .DIN(n5900),
    .DIN_t(n5900_t),
    .Q(n2203),
    .Q_t(n2203_t)
  );


  i1s3
  U4763
  (
    .DIN(n5893),
    .DIN_t(n5893_t),
    .Q(n2204),
    .Q_t(n2204_t)
  );


  i1s3
  U4764
  (
    .DIN(n5886),
    .DIN_t(n5886_t),
    .Q(n2205),
    .Q_t(n2205_t)
  );


  i1s3
  U4765
  (
    .DIN(n5879),
    .DIN_t(n5879_t),
    .Q(n2206),
    .Q_t(n2206_t)
  );


  i1s3
  U4766
  (
    .DIN(n5872),
    .DIN_t(n5872_t),
    .Q(n2207),
    .Q_t(n2207_t)
  );


  i1s3
  U4767
  (
    .DIN(n5865),
    .DIN_t(n5865_t),
    .Q(n2208),
    .Q_t(n2208_t)
  );


  i1s3
  U4768
  (
    .DIN(n6116),
    .DIN_t(n6116_t),
    .Q(n2209),
    .Q_t(n2209_t)
  );


  i1s3
  U4769
  (
    .DIN(n6117),
    .DIN_t(n6117_t),
    .Q(n2210),
    .Q_t(n2210_t)
  );


  i1s3
  U4770
  (
    .DIN(n6118),
    .DIN_t(n6118_t),
    .Q(n2211),
    .Q_t(n2211_t)
  );


  i1s3
  U4771
  (
    .DIN(n6119),
    .DIN_t(n6119_t),
    .Q(n2212),
    .Q_t(n2212_t)
  );


  i1s3
  U4772
  (
    .DIN(n6120),
    .DIN_t(n6120_t),
    .Q(n2213),
    .Q_t(n2213_t)
  );


  i1s3
  U4773
  (
    .DIN(n6121),
    .DIN_t(n6121_t),
    .Q(n2214),
    .Q_t(n2214_t)
  );


  i1s3
  U4774
  (
    .DIN(n6122),
    .DIN_t(n6122_t),
    .Q(n2215),
    .Q_t(n2215_t)
  );


  i1s3
  U4775
  (
    .DIN(n6123),
    .DIN_t(n6123_t),
    .Q(n2216),
    .Q_t(n2216_t)
  );


  i1s3
  U4776
  (
    .DIN(n6124),
    .DIN_t(n6124_t),
    .Q(n2217),
    .Q_t(n2217_t)
  );


  i1s3
  U4777
  (
    .DIN(n6125),
    .DIN_t(n6125_t),
    .Q(n2218),
    .Q_t(n2218_t)
  );


  i1s3
  U4778
  (
    .DIN(n6126),
    .DIN_t(n6126_t),
    .Q(n2219),
    .Q_t(n2219_t)
  );


  i1s3
  U4779
  (
    .DIN(n6127),
    .DIN_t(n6127_t),
    .Q(n2220),
    .Q_t(n2220_t)
  );


  i1s3
  U4780
  (
    .DIN(n6128),
    .DIN_t(n6128_t),
    .Q(n2221),
    .Q_t(n2221_t)
  );


  i1s3
  U4781
  (
    .DIN(n6129),
    .DIN_t(n6129_t),
    .Q(n2222),
    .Q_t(n2222_t)
  );


  i1s3
  U4782
  (
    .DIN(n6130),
    .DIN_t(n6130_t),
    .Q(n2223),
    .Q_t(n2223_t)
  );


  i1s3
  U4783
  (
    .DIN(n6131),
    .DIN_t(n6131_t),
    .Q(n2224),
    .Q_t(n2224_t)
  );


  i1s3
  U4784
  (
    .DIN(n6132),
    .DIN_t(n6132_t),
    .Q(n2225),
    .Q_t(n2225_t)
  );


  i1s3
  U4785
  (
    .DIN(n6133),
    .DIN_t(n6133_t),
    .Q(n2226),
    .Q_t(n2226_t)
  );


  i1s3
  U4786
  (
    .DIN(n6134),
    .DIN_t(n6134_t),
    .Q(n2227),
    .Q_t(n2227_t)
  );


  i1s3
  U4787
  (
    .DIN(n6135),
    .DIN_t(n6135_t),
    .Q(n2228),
    .Q_t(n2228_t)
  );


  i1s3
  U4788
  (
    .DIN(n6136),
    .DIN_t(n6136_t),
    .Q(n2229),
    .Q_t(n2229_t)
  );


  i1s3
  U4789
  (
    .DIN(n6137),
    .DIN_t(n6137_t),
    .Q(n2230),
    .Q_t(n2230_t)
  );


  i1s3
  U4790
  (
    .DIN(n6138),
    .DIN_t(n6138_t),
    .Q(n2231),
    .Q_t(n2231_t)
  );


  i1s3
  U4791
  (
    .DIN(n6139),
    .DIN_t(n6139_t),
    .Q(n2232),
    .Q_t(n2232_t)
  );


  i1s3
  U4792
  (
    .DIN(n6140),
    .DIN_t(n6140_t),
    .Q(n2233),
    .Q_t(n2233_t)
  );


  i1s3
  U4793
  (
    .DIN(n6141),
    .DIN_t(n6141_t),
    .Q(n2234),
    .Q_t(n2234_t)
  );


  i1s3
  U4794
  (
    .DIN(n6142),
    .DIN_t(n6142_t),
    .Q(n2235),
    .Q_t(n2235_t)
  );


  i1s3
  U4795
  (
    .DIN(n6143),
    .DIN_t(n6143_t),
    .Q(n2236),
    .Q_t(n2236_t)
  );


  i1s3
  U4796
  (
    .DIN(n6144),
    .DIN_t(n6144_t),
    .Q(n2237),
    .Q_t(n2237_t)
  );


  i1s3
  U4797
  (
    .DIN(n6145),
    .DIN_t(n6145_t),
    .Q(n2238),
    .Q_t(n2238_t)
  );


  i1s3
  U4798
  (
    .DIN(n6146),
    .DIN_t(n6146_t),
    .Q(n2239),
    .Q_t(n2239_t)
  );


  i1s3
  U4799
  (
    .DIN(n6115),
    .DIN_t(n6115_t),
    .Q(n2240),
    .Q_t(n2240_t)
  );


  i1s3
  U4800
  (
    .DIN(n6178),
    .DIN_t(n6178_t),
    .Q(n2241),
    .Q_t(n2241_t)
  );


  i1s3
  U4801
  (
    .DIN(n6147),
    .DIN_t(n6147_t),
    .Q(n2242),
    .Q_t(n2242_t)
  );


  i1s3
  U4802
  (
    .DIN(n6148),
    .DIN_t(n6148_t),
    .Q(n2243),
    .Q_t(n2243_t)
  );


  i1s3
  U4803
  (
    .DIN(n6149),
    .DIN_t(n6149_t),
    .Q(n2244),
    .Q_t(n2244_t)
  );


  i1s3
  U4804
  (
    .DIN(n6150),
    .DIN_t(n6150_t),
    .Q(n2245),
    .Q_t(n2245_t)
  );


  i1s3
  U4805
  (
    .DIN(n6151),
    .DIN_t(n6151_t),
    .Q(n2246),
    .Q_t(n2246_t)
  );


  i1s3
  U4806
  (
    .DIN(n6152),
    .DIN_t(n6152_t),
    .Q(n2247),
    .Q_t(n2247_t)
  );


  i1s3
  U4807
  (
    .DIN(n6153),
    .DIN_t(n6153_t),
    .Q(n2248),
    .Q_t(n2248_t)
  );


  i1s3
  U4808
  (
    .DIN(n6154),
    .DIN_t(n6154_t),
    .Q(n2249),
    .Q_t(n2249_t)
  );


  i1s3
  U4809
  (
    .DIN(n6155),
    .DIN_t(n6155_t),
    .Q(n2250),
    .Q_t(n2250_t)
  );


  i1s3
  U4810
  (
    .DIN(n6156),
    .DIN_t(n6156_t),
    .Q(n2251),
    .Q_t(n2251_t)
  );


  i1s3
  U4811
  (
    .DIN(n6157),
    .DIN_t(n6157_t),
    .Q(n2252),
    .Q_t(n2252_t)
  );


  i1s3
  U4812
  (
    .DIN(n6158),
    .DIN_t(n6158_t),
    .Q(n2253),
    .Q_t(n2253_t)
  );


  i1s3
  U4813
  (
    .DIN(n6159),
    .DIN_t(n6159_t),
    .Q(n2254),
    .Q_t(n2254_t)
  );


  i1s3
  U4814
  (
    .DIN(n6160),
    .DIN_t(n6160_t),
    .Q(n2255),
    .Q_t(n2255_t)
  );


  i1s3
  U4815
  (
    .DIN(n6161),
    .DIN_t(n6161_t),
    .Q(n2256),
    .Q_t(n2256_t)
  );


  i1s3
  U4816
  (
    .DIN(n6162),
    .DIN_t(n6162_t),
    .Q(n2257),
    .Q_t(n2257_t)
  );


  i1s3
  U4817
  (
    .DIN(n6163),
    .DIN_t(n6163_t),
    .Q(n2258),
    .Q_t(n2258_t)
  );


  i1s3
  U4818
  (
    .DIN(n6164),
    .DIN_t(n6164_t),
    .Q(n2259),
    .Q_t(n2259_t)
  );


  i1s3
  U4819
  (
    .DIN(n6165),
    .DIN_t(n6165_t),
    .Q(n2260),
    .Q_t(n2260_t)
  );


  i1s3
  U4820
  (
    .DIN(n6166),
    .DIN_t(n6166_t),
    .Q(n2261),
    .Q_t(n2261_t)
  );


  i1s3
  U4821
  (
    .DIN(n6167),
    .DIN_t(n6167_t),
    .Q(n2262),
    .Q_t(n2262_t)
  );


  i1s3
  U4822
  (
    .DIN(n6168),
    .DIN_t(n6168_t),
    .Q(n2263),
    .Q_t(n2263_t)
  );


  i1s3
  U4823
  (
    .DIN(n6169),
    .DIN_t(n6169_t),
    .Q(n2264),
    .Q_t(n2264_t)
  );


  i1s3
  U4824
  (
    .DIN(n6170),
    .DIN_t(n6170_t),
    .Q(n2265),
    .Q_t(n2265_t)
  );


  i1s3
  U4825
  (
    .DIN(n6171),
    .DIN_t(n6171_t),
    .Q(n2266),
    .Q_t(n2266_t)
  );


  i1s3
  U4826
  (
    .DIN(n6172),
    .DIN_t(n6172_t),
    .Q(n2267),
    .Q_t(n2267_t)
  );


  i1s3
  U4827
  (
    .DIN(n6173),
    .DIN_t(n6173_t),
    .Q(n2268),
    .Q_t(n2268_t)
  );


  i1s3
  U4828
  (
    .DIN(n6174),
    .DIN_t(n6174_t),
    .Q(n2269),
    .Q_t(n2269_t)
  );


  i1s3
  U4829
  (
    .DIN(n6175),
    .DIN_t(n6175_t),
    .Q(n2270),
    .Q_t(n2270_t)
  );


  i1s3
  U4830
  (
    .DIN(n6176),
    .DIN_t(n6176_t),
    .Q(n2271),
    .Q_t(n2271_t)
  );


  i1s3
  U4831
  (
    .DIN(n6177),
    .DIN_t(n6177_t),
    .Q(n2272),
    .Q_t(n2272_t)
  );


  i1s3
  U4832
  (
    .DIN(n6179),
    .DIN_t(n6179_t),
    .Q(n2273),
    .Q_t(n2273_t)
  );


  i1s3
  U4833
  (
    .DIN(n6180),
    .DIN_t(n6180_t),
    .Q(n2274),
    .Q_t(n2274_t)
  );


  i1s3
  U4834
  (
    .DIN(n6181),
    .DIN_t(n6181_t),
    .Q(n2275),
    .Q_t(n2275_t)
  );


  i1s3
  U4835
  (
    .DIN(n6182),
    .DIN_t(n6182_t),
    .Q(n2276),
    .Q_t(n2276_t)
  );


  i1s3
  U4836
  (
    .DIN(n6183),
    .DIN_t(n6183_t),
    .Q(n2277),
    .Q_t(n2277_t)
  );


  i1s3
  U4837
  (
    .DIN(n6184),
    .DIN_t(n6184_t),
    .Q(n2278),
    .Q_t(n2278_t)
  );


  i1s3
  U4838
  (
    .DIN(n6185),
    .DIN_t(n6185_t),
    .Q(n2279),
    .Q_t(n2279_t)
  );


  i1s3
  U4839
  (
    .DIN(n6186),
    .DIN_t(n6186_t),
    .Q(n2280),
    .Q_t(n2280_t)
  );


  i1s3
  U4840
  (
    .DIN(n6187),
    .DIN_t(n6187_t),
    .Q(n2281),
    .Q_t(n2281_t)
  );


  i1s3
  U4841
  (
    .DIN(n6188),
    .DIN_t(n6188_t),
    .Q(n2282),
    .Q_t(n2282_t)
  );


  i1s3
  U4842
  (
    .DIN(n6189),
    .DIN_t(n6189_t),
    .Q(n2283),
    .Q_t(n2283_t)
  );


  i1s3
  U4843
  (
    .DIN(n6190),
    .DIN_t(n6190_t),
    .Q(n2284),
    .Q_t(n2284_t)
  );


  i1s3
  U4844
  (
    .DIN(n6191),
    .DIN_t(n6191_t),
    .Q(n2285),
    .Q_t(n2285_t)
  );


  i1s3
  U4845
  (
    .DIN(n6192),
    .DIN_t(n6192_t),
    .Q(n2286),
    .Q_t(n2286_t)
  );


  i1s3
  U4846
  (
    .DIN(n6193),
    .DIN_t(n6193_t),
    .Q(n2287),
    .Q_t(n2287_t)
  );


  i1s3
  U4847
  (
    .DIN(n6194),
    .DIN_t(n6194_t),
    .Q(n2288),
    .Q_t(n2288_t)
  );


  i1s3
  U4848
  (
    .DIN(n6195),
    .DIN_t(n6195_t),
    .Q(n2289),
    .Q_t(n2289_t)
  );


  i1s3
  U4849
  (
    .DIN(n6196),
    .DIN_t(n6196_t),
    .Q(n2290),
    .Q_t(n2290_t)
  );


  i1s3
  U4850
  (
    .DIN(n6286),
    .DIN_t(n6286_t),
    .Q(n2291),
    .Q_t(n2291_t)
  );


  i1s3
  U4851
  (
    .DIN(n6342),
    .DIN_t(n6342_t),
    .Q(n2292),
    .Q_t(n2292_t)
  );


  i1s3
  U4852
  (
    .DIN(n6354),
    .DIN_t(n6354_t),
    .Q(n2293),
    .Q_t(n2293_t)
  );


  i1s3
  U4853
  (
    .DIN(n6376),
    .DIN_t(n6376_t),
    .Q(n2294),
    .Q_t(n2294_t)
  );


  i1s3
  U4854
  (
    .DIN(n6377),
    .DIN_t(n6377_t),
    .Q(n2295),
    .Q_t(n2295_t)
  );


  i1s3
  U4855
  (
    .DIN(n6378),
    .DIN_t(n6378_t),
    .Q(n2296),
    .Q_t(n2296_t)
  );


  i1s3
  U4856
  (
    .DIN(n6379),
    .DIN_t(n6379_t),
    .Q(n2297),
    .Q_t(n2297_t)
  );


  i1s3
  U4857
  (
    .DIN(n6380),
    .DIN_t(n6380_t),
    .Q(n2298),
    .Q_t(n2298_t)
  );


  i1s3
  U4858
  (
    .DIN(n6381),
    .DIN_t(n6381_t),
    .Q(n2299),
    .Q_t(n2299_t)
  );


  i1s3
  U4859
  (
    .DIN(n6382),
    .DIN_t(n6382_t),
    .Q(n2300),
    .Q_t(n2300_t)
  );


  i1s3
  U4860
  (
    .DIN(n6431),
    .DIN_t(n6431_t),
    .Q(n2301),
    .Q_t(n2301_t)
  );


  i1s3
  U4861
  (
    .DIN(n6432),
    .DIN_t(n6432_t),
    .Q(n2302),
    .Q_t(n2302_t)
  );


  i1s3
  U4862
  (
    .DIN(n6433),
    .DIN_t(n6433_t),
    .Q(n2303),
    .Q_t(n2303_t)
  );


  i1s3
  U4863
  (
    .DIN(n6434),
    .DIN_t(n6434_t),
    .Q(n2304),
    .Q_t(n2304_t)
  );


  i1s3
  U4866
  (
    .DIN(TM1),
    .DIN_t(TM1_t),
    .Q(n2307),
    .Q_t(n2307_t)
  );


  ib1s9
  U4867
  (
    .DIN(n6593),
    .DIN_t(n6593_t),
    .Q(n6563),
    .Q_t(n6563_t)
  );


  ib1s9
  U4868
  (
    .DIN(n6593),
    .DIN_t(n6593_t),
    .Q(n6564),
    .Q_t(n6564_t)
  );


  ib1s9
  U4869
  (
    .DIN(n6592),
    .DIN_t(n6592_t),
    .Q(n6565),
    .Q_t(n6565_t)
  );


  ib1s9
  U4870
  (
    .DIN(n6592),
    .DIN_t(n6592_t),
    .Q(n6566),
    .Q_t(n6566_t)
  );


  ib1s9
  U4871
  (
    .DIN(n6592),
    .DIN_t(n6592_t),
    .Q(n6567),
    .Q_t(n6567_t)
  );


  ib1s9
  U4872
  (
    .DIN(n6591),
    .DIN_t(n6591_t),
    .Q(n6568),
    .Q_t(n6568_t)
  );


  ib1s9
  U4873
  (
    .DIN(n6591),
    .DIN_t(n6591_t),
    .Q(n6569),
    .Q_t(n6569_t)
  );


  ib1s9
  U4874
  (
    .DIN(n6591),
    .DIN_t(n6591_t),
    .Q(n6570),
    .Q_t(n6570_t)
  );


  ib1s9
  U4875
  (
    .DIN(n6590),
    .DIN_t(n6590_t),
    .Q(n6571),
    .Q_t(n6571_t)
  );


  ib1s9
  U4876
  (
    .DIN(n6590),
    .DIN_t(n6590_t),
    .Q(n6572),
    .Q_t(n6572_t)
  );


  ib1s9
  U4877
  (
    .DIN(n6590),
    .DIN_t(n6590_t),
    .Q(n6573),
    .Q_t(n6573_t)
  );


  ib1s9
  U4878
  (
    .DIN(n6589),
    .DIN_t(n6589_t),
    .Q(n6574),
    .Q_t(n6574_t)
  );


  ib1s9
  U4879
  (
    .DIN(n6589),
    .DIN_t(n6589_t),
    .Q(n6575),
    .Q_t(n6575_t)
  );


  ib1s9
  U4880
  (
    .DIN(n6589),
    .DIN_t(n6589_t),
    .Q(n6576),
    .Q_t(n6576_t)
  );


  ib1s9
  U4881
  (
    .DIN(n6588),
    .DIN_t(n6588_t),
    .Q(n6577),
    .Q_t(n6577_t)
  );


  ib1s9
  U4882
  (
    .DIN(n6588),
    .DIN_t(n6588_t),
    .Q(n6578),
    .Q_t(n6578_t)
  );


  ib1s9
  U4883
  (
    .DIN(n6588),
    .DIN_t(n6588_t),
    .Q(n6579),
    .Q_t(n6579_t)
  );


  ib1s9
  U4884
  (
    .DIN(n6587),
    .DIN_t(n6587_t),
    .Q(n6580),
    .Q_t(n6580_t)
  );


  ib1s9
  U4885
  (
    .DIN(n6587),
    .DIN_t(n6587_t),
    .Q(n6581),
    .Q_t(n6581_t)
  );


  ib1s9
  U4886
  (
    .DIN(n6587),
    .DIN_t(n6587_t),
    .Q(n6582),
    .Q_t(n6582_t)
  );


  ib1s9
  U4887
  (
    .DIN(n6586),
    .DIN_t(n6586_t),
    .Q(n6583),
    .Q_t(n6583_t)
  );


  ib1s9
  U4888
  (
    .DIN(n6586),
    .DIN_t(n6586_t),
    .Q(n6584),
    .Q_t(n6584_t)
  );


  ib1s9
  U4889
  (
    .DIN(n6624),
    .DIN_t(n6624_t),
    .Q(n6594),
    .Q_t(n6594_t)
  );


  ib1s9
  U4890
  (
    .DIN(n6624),
    .DIN_t(n6624_t),
    .Q(n6595),
    .Q_t(n6595_t)
  );


  ib1s9
  U4891
  (
    .DIN(n6623),
    .DIN_t(n6623_t),
    .Q(n6596),
    .Q_t(n6596_t)
  );


  ib1s9
  U4892
  (
    .DIN(n6623),
    .DIN_t(n6623_t),
    .Q(n6597),
    .Q_t(n6597_t)
  );


  ib1s9
  U4893
  (
    .DIN(n6623),
    .DIN_t(n6623_t),
    .Q(n6598),
    .Q_t(n6598_t)
  );


  ib1s9
  U4894
  (
    .DIN(n6622),
    .DIN_t(n6622_t),
    .Q(n6599),
    .Q_t(n6599_t)
  );


  ib1s9
  U4895
  (
    .DIN(n6622),
    .DIN_t(n6622_t),
    .Q(n6600),
    .Q_t(n6600_t)
  );


  ib1s9
  U4896
  (
    .DIN(n6622),
    .DIN_t(n6622_t),
    .Q(n6601),
    .Q_t(n6601_t)
  );


  ib1s9
  U4897
  (
    .DIN(n6621),
    .DIN_t(n6621_t),
    .Q(n6602),
    .Q_t(n6602_t)
  );


  ib1s9
  U4898
  (
    .DIN(n6621),
    .DIN_t(n6621_t),
    .Q(n6603),
    .Q_t(n6603_t)
  );


  ib1s9
  U4899
  (
    .DIN(n6621),
    .DIN_t(n6621_t),
    .Q(n6604),
    .Q_t(n6604_t)
  );


  ib1s9
  U4900
  (
    .DIN(n6620),
    .DIN_t(n6620_t),
    .Q(n6605),
    .Q_t(n6605_t)
  );


  ib1s9
  U4901
  (
    .DIN(n6620),
    .DIN_t(n6620_t),
    .Q(n6606),
    .Q_t(n6606_t)
  );


  ib1s9
  U4902
  (
    .DIN(n6620),
    .DIN_t(n6620_t),
    .Q(n6607),
    .Q_t(n6607_t)
  );


  ib1s9
  U4903
  (
    .DIN(n6619),
    .DIN_t(n6619_t),
    .Q(n6608),
    .Q_t(n6608_t)
  );


  ib1s9
  U4904
  (
    .DIN(n6619),
    .DIN_t(n6619_t),
    .Q(n6609),
    .Q_t(n6609_t)
  );


  ib1s9
  U4905
  (
    .DIN(n6619),
    .DIN_t(n6619_t),
    .Q(n6610),
    .Q_t(n6610_t)
  );


  ib1s9
  U4906
  (
    .DIN(n6618),
    .DIN_t(n6618_t),
    .Q(n6611),
    .Q_t(n6611_t)
  );


  ib1s9
  U4907
  (
    .DIN(n6618),
    .DIN_t(n6618_t),
    .Q(n6612),
    .Q_t(n6612_t)
  );


  ib1s9
  U4908
  (
    .DIN(n6618),
    .DIN_t(n6618_t),
    .Q(n6613),
    .Q_t(n6613_t)
  );


  ib1s9
  U4909
  (
    .DIN(n6617),
    .DIN_t(n6617_t),
    .Q(n6614),
    .Q_t(n6614_t)
  );


  ib1s9
  U4910
  (
    .DIN(n6617),
    .DIN_t(n6617_t),
    .Q(n6615),
    .Q_t(n6615_t)
  );


  ib1s9
  U4911
  (
    .DIN(n6655),
    .DIN_t(n6655_t),
    .Q(n6625),
    .Q_t(n6625_t)
  );


  ib1s9
  U4912
  (
    .DIN(n6655),
    .DIN_t(n6655_t),
    .Q(n6626),
    .Q_t(n6626_t)
  );


  ib1s9
  U4913
  (
    .DIN(n6654),
    .DIN_t(n6654_t),
    .Q(n6627),
    .Q_t(n6627_t)
  );


  ib1s9
  U4914
  (
    .DIN(n6654),
    .DIN_t(n6654_t),
    .Q(n6628),
    .Q_t(n6628_t)
  );


  ib1s9
  U4915
  (
    .DIN(n6654),
    .DIN_t(n6654_t),
    .Q(n6629),
    .Q_t(n6629_t)
  );


  ib1s9
  U4916
  (
    .DIN(n6653),
    .DIN_t(n6653_t),
    .Q(n6630),
    .Q_t(n6630_t)
  );


  ib1s9
  U4917
  (
    .DIN(n6653),
    .DIN_t(n6653_t),
    .Q(n6631),
    .Q_t(n6631_t)
  );


  ib1s9
  U4918
  (
    .DIN(n6653),
    .DIN_t(n6653_t),
    .Q(n6632),
    .Q_t(n6632_t)
  );


  ib1s9
  U4919
  (
    .DIN(n6652),
    .DIN_t(n6652_t),
    .Q(n6633),
    .Q_t(n6633_t)
  );


  ib1s9
  U4920
  (
    .DIN(n6652),
    .DIN_t(n6652_t),
    .Q(n6634),
    .Q_t(n6634_t)
  );


  ib1s9
  U4921
  (
    .DIN(n6652),
    .DIN_t(n6652_t),
    .Q(n6635),
    .Q_t(n6635_t)
  );


  ib1s9
  U4922
  (
    .DIN(n6651),
    .DIN_t(n6651_t),
    .Q(n6636),
    .Q_t(n6636_t)
  );


  ib1s9
  U4923
  (
    .DIN(n6651),
    .DIN_t(n6651_t),
    .Q(n6637),
    .Q_t(n6637_t)
  );


  ib1s9
  U4924
  (
    .DIN(n6651),
    .DIN_t(n6651_t),
    .Q(n6638),
    .Q_t(n6638_t)
  );


  ib1s9
  U4925
  (
    .DIN(n6650),
    .DIN_t(n6650_t),
    .Q(n6639),
    .Q_t(n6639_t)
  );


  ib1s9
  U4926
  (
    .DIN(n6650),
    .DIN_t(n6650_t),
    .Q(n6640),
    .Q_t(n6640_t)
  );


  ib1s9
  U4927
  (
    .DIN(n6650),
    .DIN_t(n6650_t),
    .Q(n6641),
    .Q_t(n6641_t)
  );


  ib1s9
  U4928
  (
    .DIN(n6649),
    .DIN_t(n6649_t),
    .Q(n6642),
    .Q_t(n6642_t)
  );


  ib1s9
  U4929
  (
    .DIN(n6649),
    .DIN_t(n6649_t),
    .Q(n6643),
    .Q_t(n6643_t)
  );


  ib1s9
  U4930
  (
    .DIN(n6649),
    .DIN_t(n6649_t),
    .Q(n6644),
    .Q_t(n6644_t)
  );


  ib1s9
  U4931
  (
    .DIN(n6648),
    .DIN_t(n6648_t),
    .Q(n6645),
    .Q_t(n6645_t)
  );


  ib1s9
  U4932
  (
    .DIN(n6648),
    .DIN_t(n6648_t),
    .Q(n6646),
    .Q_t(n6646_t)
  );


  ib1s9
  U4933
  (
    .DIN(n6686),
    .DIN_t(n6686_t),
    .Q(n6656),
    .Q_t(n6656_t)
  );


  ib1s9
  U4934
  (
    .DIN(n6686),
    .DIN_t(n6686_t),
    .Q(n6657),
    .Q_t(n6657_t)
  );


  ib1s9
  U4935
  (
    .DIN(n6685),
    .DIN_t(n6685_t),
    .Q(n6658),
    .Q_t(n6658_t)
  );


  ib1s9
  U4936
  (
    .DIN(n6685),
    .DIN_t(n6685_t),
    .Q(n6659),
    .Q_t(n6659_t)
  );


  ib1s9
  U4937
  (
    .DIN(n6685),
    .DIN_t(n6685_t),
    .Q(n6660),
    .Q_t(n6660_t)
  );


  ib1s9
  U4938
  (
    .DIN(n6684),
    .DIN_t(n6684_t),
    .Q(n6661),
    .Q_t(n6661_t)
  );


  ib1s9
  U4939
  (
    .DIN(n6684),
    .DIN_t(n6684_t),
    .Q(n6662),
    .Q_t(n6662_t)
  );


  ib1s9
  U4940
  (
    .DIN(n6684),
    .DIN_t(n6684_t),
    .Q(n6663),
    .Q_t(n6663_t)
  );


  ib1s9
  U4941
  (
    .DIN(n6683),
    .DIN_t(n6683_t),
    .Q(n6664),
    .Q_t(n6664_t)
  );


  ib1s9
  U4942
  (
    .DIN(n6683),
    .DIN_t(n6683_t),
    .Q(n6665),
    .Q_t(n6665_t)
  );


  ib1s9
  U4943
  (
    .DIN(n6683),
    .DIN_t(n6683_t),
    .Q(n6666),
    .Q_t(n6666_t)
  );


  ib1s9
  U4944
  (
    .DIN(n6682),
    .DIN_t(n6682_t),
    .Q(n6667),
    .Q_t(n6667_t)
  );


  ib1s9
  U4945
  (
    .DIN(n6682),
    .DIN_t(n6682_t),
    .Q(n6668),
    .Q_t(n6668_t)
  );


  ib1s9
  U4946
  (
    .DIN(n6682),
    .DIN_t(n6682_t),
    .Q(n6669),
    .Q_t(n6669_t)
  );


  ib1s9
  U4947
  (
    .DIN(n6681),
    .DIN_t(n6681_t),
    .Q(n6670),
    .Q_t(n6670_t)
  );


  ib1s9
  U4948
  (
    .DIN(n6681),
    .DIN_t(n6681_t),
    .Q(n6671),
    .Q_t(n6671_t)
  );


  ib1s9
  U4949
  (
    .DIN(n6681),
    .DIN_t(n6681_t),
    .Q(n6672),
    .Q_t(n6672_t)
  );


  ib1s9
  U4950
  (
    .DIN(n6680),
    .DIN_t(n6680_t),
    .Q(n6673),
    .Q_t(n6673_t)
  );


  ib1s9
  U4951
  (
    .DIN(n6680),
    .DIN_t(n6680_t),
    .Q(n6674),
    .Q_t(n6674_t)
  );


  ib1s9
  U4952
  (
    .DIN(n6680),
    .DIN_t(n6680_t),
    .Q(n6675),
    .Q_t(n6675_t)
  );


  ib1s9
  U4953
  (
    .DIN(n6679),
    .DIN_t(n6679_t),
    .Q(n6676),
    .Q_t(n6676_t)
  );


  ib1s9
  U4954
  (
    .DIN(n6679),
    .DIN_t(n6679_t),
    .Q(n6677),
    .Q_t(n6677_t)
  );


  ib1s9
  U4955
  (
    .DIN(n6702),
    .DIN_t(n6702_t),
    .Q(n6687),
    .Q_t(n6687_t)
  );


  ib1s9
  U4956
  (
    .DIN(n6702),
    .DIN_t(n6702_t),
    .Q(n6688),
    .Q_t(n6688_t)
  );


  ib1s9
  U4957
  (
    .DIN(n6702),
    .DIN_t(n6702_t),
    .Q(n6689),
    .Q_t(n6689_t)
  );


  ib1s9
  U4958
  (
    .DIN(n6701),
    .DIN_t(n6701_t),
    .Q(n6690),
    .Q_t(n6690_t)
  );


  ib1s9
  U4959
  (
    .DIN(n6701),
    .DIN_t(n6701_t),
    .Q(n6691),
    .Q_t(n6691_t)
  );


  ib1s9
  U4960
  (
    .DIN(n6701),
    .DIN_t(n6701_t),
    .Q(n6692),
    .Q_t(n6692_t)
  );


  ib1s9
  U4961
  (
    .DIN(n6700),
    .DIN_t(n6700_t),
    .Q(n6693),
    .Q_t(n6693_t)
  );


  ib1s9
  U4962
  (
    .DIN(n6700),
    .DIN_t(n6700_t),
    .Q(n6694),
    .Q_t(n6694_t)
  );


  ib1s9
  U4963
  (
    .DIN(n6700),
    .DIN_t(n6700_t),
    .Q(n6695),
    .Q_t(n6695_t)
  );


  ib1s9
  U4964
  (
    .DIN(n6699),
    .DIN_t(n6699_t),
    .Q(n6696),
    .Q_t(n6696_t)
  );


  ib1s9
  U4965
  (
    .DIN(n6699),
    .DIN_t(n6699_t),
    .Q(n6697),
    .Q_t(n6697_t)
  );


  ib1s9
  U4966
  (
    .DIN(n6706),
    .DIN_t(n6706_t),
    .Q(n6703),
    .Q_t(n6703_t)
  );


  ib1s9
  U4967
  (
    .DIN(n6706),
    .DIN_t(n6706_t),
    .Q(n6704),
    .Q_t(n6704_t)
  );


  ib1s9
  U4968
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6712),
    .Q_t(n6712_t)
  );


  ib1s9
  U4969
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6713),
    .Q_t(n6713_t)
  );


  ib1s9
  U4970
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6714),
    .Q_t(n6714_t)
  );


  ib1s9
  U4971
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6715),
    .Q_t(n6715_t)
  );


  ib1s9
  U4972
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6716),
    .Q_t(n6716_t)
  );


  ib1s9
  U4973
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6717),
    .Q_t(n6717_t)
  );


  ib1s9
  U4974
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6718),
    .Q_t(n6718_t)
  );


  ib1s9
  U4975
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6719),
    .Q_t(n6719_t)
  );


  ib1s9
  U4976
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6720),
    .Q_t(n6720_t)
  );


  ib1s9
  U4977
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6721),
    .Q_t(n6721_t)
  );


  ib1s9
  U4978
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6722),
    .Q_t(n6722_t)
  );


  ib1s9
  U4979
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6723),
    .Q_t(n6723_t)
  );


  ib1s9
  U4980
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6724),
    .Q_t(n6724_t)
  );


  ib1s9
  U4981
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6725),
    .Q_t(n6725_t)
  );


  ib1s9
  U4982
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6726),
    .Q_t(n6726_t)
  );


  ib1s9
  U4983
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6727),
    .Q_t(n6727_t)
  );


  ib1s9
  U4984
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6728),
    .Q_t(n6728_t)
  );


  ib1s9
  U4985
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6729),
    .Q_t(n6729_t)
  );


  ib1s9
  U4986
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6730),
    .Q_t(n6730_t)
  );


  ib1s9
  U4987
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6731),
    .Q_t(n6731_t)
  );


  ib1s9
  U4988
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6732),
    .Q_t(n6732_t)
  );


  ib1s9
  U4989
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6733),
    .Q_t(n6733_t)
  );


  ib1s9
  U4990
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6734),
    .Q_t(n6734_t)
  );


  ib1s9
  U4991
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6735),
    .Q_t(n6735_t)
  );


  ib1s9
  U4992
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6736),
    .Q_t(n6736_t)
  );


  ib1s9
  U4993
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6737),
    .Q_t(n6737_t)
  );


  ib1s9
  U4994
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6738),
    .Q_t(n6738_t)
  );


  ib1s9
  U4995
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6739),
    .Q_t(n6739_t)
  );


  ib1s9
  U4996
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6740),
    .Q_t(n6740_t)
  );


  ib1s9
  U4997
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6741),
    .Q_t(n6741_t)
  );


  ib1s9
  U4998
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6742),
    .Q_t(n6742_t)
  );


  ib1s9
  U4999
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6743),
    .Q_t(n6743_t)
  );


  ib1s9
  U5000
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6744),
    .Q_t(n6744_t)
  );


  ib1s9
  U5001
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6745),
    .Q_t(n6745_t)
  );


  ib1s9
  U5002
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6746),
    .Q_t(n6746_t)
  );


  ib1s9
  U5003
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6747),
    .Q_t(n6747_t)
  );


  ib1s9
  U5004
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6748),
    .Q_t(n6748_t)
  );


  ib1s9
  U5005
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6749),
    .Q_t(n6749_t)
  );


  ib1s9
  U5006
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6750),
    .Q_t(n6750_t)
  );


  ib1s9
  U5007
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6751),
    .Q_t(n6751_t)
  );


  ib1s9
  U5008
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6752),
    .Q_t(n6752_t)
  );


  ib1s9
  U5009
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6753),
    .Q_t(n6753_t)
  );


  ib1s9
  U5010
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6754),
    .Q_t(n6754_t)
  );


  ib1s9
  U5011
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6755),
    .Q_t(n6755_t)
  );


  ib1s9
  U5012
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6756),
    .Q_t(n6756_t)
  );


  ib1s9
  U5013
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6757),
    .Q_t(n6757_t)
  );


  ib1s9
  U5014
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6758),
    .Q_t(n6758_t)
  );


  ib1s9
  U5015
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6759),
    .Q_t(n6759_t)
  );


  ib1s9
  U5016
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6760),
    .Q_t(n6760_t)
  );


  ib1s9
  U5017
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6761),
    .Q_t(n6761_t)
  );


  ib1s9
  U5018
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6762),
    .Q_t(n6762_t)
  );


  ib1s9
  U5019
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6763),
    .Q_t(n6763_t)
  );


  ib1s9
  U5020
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6764),
    .Q_t(n6764_t)
  );


  ib1s9
  U5021
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6765),
    .Q_t(n6765_t)
  );


  ib1s9
  U5022
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6766),
    .Q_t(n6766_t)
  );


  ib1s9
  U5023
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6767),
    .Q_t(n6767_t)
  );


  ib1s9
  U5024
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6768),
    .Q_t(n6768_t)
  );


  ib1s9
  U5025
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6769),
    .Q_t(n6769_t)
  );


  ib1s9
  U5026
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6770),
    .Q_t(n6770_t)
  );


  ib1s9
  U5027
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6771),
    .Q_t(n6771_t)
  );


  ib1s9
  U5028
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6772),
    .Q_t(n6772_t)
  );


  ib1s9
  U5029
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6773),
    .Q_t(n6773_t)
  );


  ib1s9
  U5030
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6774),
    .Q_t(n6774_t)
  );


  ib1s9
  U5031
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6775),
    .Q_t(n6775_t)
  );


  ib1s9
  U5032
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6776),
    .Q_t(n6776_t)
  );


  ib1s9
  U5033
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6777),
    .Q_t(n6777_t)
  );


  ib1s9
  U5034
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6778),
    .Q_t(n6778_t)
  );


  ib1s9
  U5035
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6779),
    .Q_t(n6779_t)
  );


  ib1s9
  U5036
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6780),
    .Q_t(n6780_t)
  );


  ib1s9
  U5037
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6781),
    .Q_t(n6781_t)
  );


  ib1s9
  U5038
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6782),
    .Q_t(n6782_t)
  );


  ib1s9
  U5039
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6783),
    .Q_t(n6783_t)
  );


  ib1s9
  U5040
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6784),
    .Q_t(n6784_t)
  );


  ib1s9
  U5041
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6785),
    .Q_t(n6785_t)
  );


  ib1s9
  U5042
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6786),
    .Q_t(n6786_t)
  );


  ib1s9
  U5043
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6787),
    .Q_t(n6787_t)
  );


  ib1s9
  U5044
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6788),
    .Q_t(n6788_t)
  );


  ib1s9
  U5045
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6789),
    .Q_t(n6789_t)
  );


  ib1s9
  U5046
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6790),
    .Q_t(n6790_t)
  );


  ib1s9
  U5047
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6791),
    .Q_t(n6791_t)
  );


  ib1s9
  U5048
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6792),
    .Q_t(n6792_t)
  );


  ib1s9
  U5049
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6793),
    .Q_t(n6793_t)
  );


  ib1s9
  U5050
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6794),
    .Q_t(n6794_t)
  );


  ib1s9
  U5051
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6795),
    .Q_t(n6795_t)
  );


  ib1s9
  U5052
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6796),
    .Q_t(n6796_t)
  );


  ib1s9
  U5053
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6797),
    .Q_t(n6797_t)
  );


  ib1s9
  U5054
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6798),
    .Q_t(n6798_t)
  );


  ib1s9
  U5055
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6799),
    .Q_t(n6799_t)
  );


  ib1s9
  U5056
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6800),
    .Q_t(n6800_t)
  );


  ib1s9
  U5057
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6801),
    .Q_t(n6801_t)
  );


  ib1s9
  U5058
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6802),
    .Q_t(n6802_t)
  );


  ib1s9
  U5059
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6803),
    .Q_t(n6803_t)
  );


  ib1s9
  U5060
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6804),
    .Q_t(n6804_t)
  );


  ib1s9
  U5061
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6805),
    .Q_t(n6805_t)
  );


  ib1s9
  U5062
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6806),
    .Q_t(n6806_t)
  );


  ib1s9
  U5063
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6807),
    .Q_t(n6807_t)
  );


  ib1s9
  U5064
  (
    .DIN(RESET),
    .DIN_t(RESET_t),
    .Q(n6808),
    .Q_t(n6808_t)
  );


  i1s11
  U5065
  (
    .DIN(n6586),
    .DIN_t(n6586_t),
    .Q(n6585),
    .Q_t(n6585_t)
  );


  i1s11
  U5066
  (
    .DIN(n2317),
    .DIN_t(n2317_t),
    .Q(n6586),
    .Q_t(n6586_t)
  );


  i1s11
  U5067
  (
    .DIN(n2317),
    .DIN_t(n2317_t),
    .Q(n6587),
    .Q_t(n6587_t)
  );


  i1s11
  U5068
  (
    .DIN(n2317),
    .DIN_t(n2317_t),
    .Q(n6588),
    .Q_t(n6588_t)
  );


  i1s11
  U5069
  (
    .DIN(n2317),
    .DIN_t(n2317_t),
    .Q(n6589),
    .Q_t(n6589_t)
  );


  i1s11
  U5070
  (
    .DIN(n2317),
    .DIN_t(n2317_t),
    .Q(n6590),
    .Q_t(n6590_t)
  );


  i1s11
  U5071
  (
    .DIN(n2317),
    .DIN_t(n2317_t),
    .Q(n6591),
    .Q_t(n6591_t)
  );


  i1s11
  U5072
  (
    .DIN(n2317),
    .DIN_t(n2317_t),
    .Q(n6592),
    .Q_t(n6592_t)
  );


  i1s11
  U5073
  (
    .DIN(n2317),
    .DIN_t(n2317_t),
    .Q(n6593),
    .Q_t(n6593_t)
  );


  i1s11
  U5074
  (
    .DIN(n6617),
    .DIN_t(n6617_t),
    .Q(n6616),
    .Q_t(n6616_t)
  );


  i1s11
  U5075
  (
    .DIN(n2316),
    .DIN_t(n2316_t),
    .Q(n6617),
    .Q_t(n6617_t)
  );


  i1s11
  U5076
  (
    .DIN(n2316),
    .DIN_t(n2316_t),
    .Q(n6618),
    .Q_t(n6618_t)
  );


  i1s11
  U5077
  (
    .DIN(n2316),
    .DIN_t(n2316_t),
    .Q(n6619),
    .Q_t(n6619_t)
  );


  i1s11
  U5078
  (
    .DIN(n2316),
    .DIN_t(n2316_t),
    .Q(n6620),
    .Q_t(n6620_t)
  );


  i1s11
  U5079
  (
    .DIN(n2316),
    .DIN_t(n2316_t),
    .Q(n6621),
    .Q_t(n6621_t)
  );


  i1s11
  U5080
  (
    .DIN(n2316),
    .DIN_t(n2316_t),
    .Q(n6622),
    .Q_t(n6622_t)
  );


  i1s11
  U5081
  (
    .DIN(n2316),
    .DIN_t(n2316_t),
    .Q(n6623),
    .Q_t(n6623_t)
  );


  i1s11
  U5082
  (
    .DIN(n2316),
    .DIN_t(n2316_t),
    .Q(n6624),
    .Q_t(n6624_t)
  );


  i1s11
  U5083
  (
    .DIN(n6648),
    .DIN_t(n6648_t),
    .Q(n6647),
    .Q_t(n6647_t)
  );


  i1s11
  U5084
  (
    .DIN(n2314),
    .DIN_t(n2314_t),
    .Q(n6648),
    .Q_t(n6648_t)
  );


  i1s11
  U5085
  (
    .DIN(n2314),
    .DIN_t(n2314_t),
    .Q(n6649),
    .Q_t(n6649_t)
  );


  i1s11
  U5086
  (
    .DIN(n2314),
    .DIN_t(n2314_t),
    .Q(n6650),
    .Q_t(n6650_t)
  );


  i1s11
  U5087
  (
    .DIN(n2314),
    .DIN_t(n2314_t),
    .Q(n6651),
    .Q_t(n6651_t)
  );


  i1s11
  U5088
  (
    .DIN(n2314),
    .DIN_t(n2314_t),
    .Q(n6652),
    .Q_t(n6652_t)
  );


  i1s11
  U5089
  (
    .DIN(n2314),
    .DIN_t(n2314_t),
    .Q(n6653),
    .Q_t(n6653_t)
  );


  i1s11
  U5090
  (
    .DIN(n2314),
    .DIN_t(n2314_t),
    .Q(n6654),
    .Q_t(n6654_t)
  );


  i1s11
  U5091
  (
    .DIN(n2314),
    .DIN_t(n2314_t),
    .Q(n6655),
    .Q_t(n6655_t)
  );


  i1s11
  U5092
  (
    .DIN(n6679),
    .DIN_t(n6679_t),
    .Q(n6678),
    .Q_t(n6678_t)
  );


  i1s11
  U5093
  (
    .DIN(n2312),
    .DIN_t(n2312_t),
    .Q(n6679),
    .Q_t(n6679_t)
  );


  i1s11
  U5094
  (
    .DIN(n2312),
    .DIN_t(n2312_t),
    .Q(n6680),
    .Q_t(n6680_t)
  );


  i1s11
  U5095
  (
    .DIN(n2312),
    .DIN_t(n2312_t),
    .Q(n6681),
    .Q_t(n6681_t)
  );


  i1s11
  U5096
  (
    .DIN(n2312),
    .DIN_t(n2312_t),
    .Q(n6682),
    .Q_t(n6682_t)
  );


  i1s11
  U5097
  (
    .DIN(n2312),
    .DIN_t(n2312_t),
    .Q(n6683),
    .Q_t(n6683_t)
  );


  i1s11
  U5098
  (
    .DIN(n2312),
    .DIN_t(n2312_t),
    .Q(n6684),
    .Q_t(n6684_t)
  );


  i1s11
  U5099
  (
    .DIN(n2312),
    .DIN_t(n2312_t),
    .Q(n6685),
    .Q_t(n6685_t)
  );


  i1s11
  U5100
  (
    .DIN(n2312),
    .DIN_t(n2312_t),
    .Q(n6686),
    .Q_t(n6686_t)
  );


  i1s12
  U5101
  (
    .DIN(n6699),
    .DIN_t(n6699_t),
    .Q(n6698),
    .Q_t(n6698_t)
  );


  i1s12
  U5102
  (
    .DIN(n2307),
    .DIN_t(n2307_t),
    .Q(n6699),
    .Q_t(n6699_t)
  );


  i1s12
  U5103
  (
    .DIN(n2307),
    .DIN_t(n2307_t),
    .Q(n6700),
    .Q_t(n6700_t)
  );


  i1s12
  U5104
  (
    .DIN(n2307),
    .DIN_t(n2307_t),
    .Q(n6701),
    .Q_t(n6701_t)
  );


  i1s12
  U5105
  (
    .DIN(n2307),
    .DIN_t(n2307_t),
    .Q(n6702),
    .Q_t(n6702_t)
  );


  i1s12
  U5106
  (
    .DIN(n6706),
    .DIN_t(n6706_t),
    .Q(n6705),
    .Q_t(n6705_t)
  );


  i1s12
  U5107
  (
    .DIN(TM0),
    .DIN_t(TM0_t),
    .Q(n6706),
    .Q_t(n6706_t)
  );


  i1s12
  U5108
  (
    .DIN(TM0),
    .DIN_t(TM0_t),
    .Q(n6707),
    .Q_t(n6707_t)
  );


  i1s12
  U5109
  (
    .DIN(TM0),
    .DIN_t(TM0_t),
    .Q(n6708),
    .Q_t(n6708_t)
  );


  i1s12
  U5110
  (
    .DIN(TM0),
    .DIN_t(TM0_t),
    .Q(n6709),
    .Q_t(n6709_t)
  );


  i1s12
  U5111
  (
    .DIN(TM0),
    .DIN_t(TM0_t),
    .Q(n6710),
    .Q_t(n6710_t)
  );


  i1s12
  U5112
  (
    .DIN(TM0),
    .DIN_t(TM0_t),
    .Q(n6711),
    .Q_t(n6711_t)
  );


  sdffs1
  \DFF_1727/Q_reg 
  (
    .DIN(WX11670),
    .DIN_t(WX11670_t),
    .SDIN(CRC_OUT_1_30),
    .SDIN_t(CRC_OUT_1_30_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_31),
    .Q_t(CRC_OUT_1_31_t),
    .QN(n6337),
    .QN_t(n6337_t)
  );


  sdffs1
  \DFF_1726/Q_reg 
  (
    .DIN(WX11668),
    .DIN_t(WX11668_t),
    .SDIN(CRC_OUT_1_29),
    .SDIN_t(CRC_OUT_1_29_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_30),
    .Q_t(CRC_OUT_1_30_t),
    .QN(n6336),
    .QN_t(n6336_t)
  );


  sdffs1
  \DFF_1725/Q_reg 
  (
    .DIN(WX11666),
    .DIN_t(WX11666_t),
    .SDIN(CRC_OUT_1_28),
    .SDIN_t(CRC_OUT_1_28_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_29),
    .Q_t(CRC_OUT_1_29_t),
    .QN(n6331),
    .QN_t(n6331_t)
  );


  sdffs1
  \DFF_1724/Q_reg 
  (
    .DIN(WX11664),
    .DIN_t(WX11664_t),
    .SDIN(CRC_OUT_1_27),
    .SDIN_t(CRC_OUT_1_27_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_28),
    .Q_t(CRC_OUT_1_28_t),
    .QN(n6326),
    .QN_t(n6326_t)
  );


  sdffs1
  \DFF_1723/Q_reg 
  (
    .DIN(WX11662),
    .DIN_t(WX11662_t),
    .SDIN(CRC_OUT_1_26),
    .SDIN_t(CRC_OUT_1_26_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_27),
    .Q_t(CRC_OUT_1_27_t),
    .QN(n6321),
    .QN_t(n6321_t)
  );


  sdffs1
  \DFF_1722/Q_reg 
  (
    .DIN(WX11660),
    .DIN_t(WX11660_t),
    .SDIN(CRC_OUT_1_25),
    .SDIN_t(CRC_OUT_1_25_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_26),
    .Q_t(CRC_OUT_1_26_t),
    .QN(n6316),
    .QN_t(n6316_t)
  );


  sdffs1
  \DFF_1721/Q_reg 
  (
    .DIN(WX11658),
    .DIN_t(WX11658_t),
    .SDIN(CRC_OUT_1_24),
    .SDIN_t(CRC_OUT_1_24_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_25),
    .Q_t(CRC_OUT_1_25_t),
    .QN(n6311),
    .QN_t(n6311_t)
  );


  sdffs1
  \DFF_1720/Q_reg 
  (
    .DIN(WX11656),
    .DIN_t(WX11656_t),
    .SDIN(CRC_OUT_1_23),
    .SDIN_t(CRC_OUT_1_23_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_24),
    .Q_t(CRC_OUT_1_24_t),
    .QN(n6306),
    .QN_t(n6306_t)
  );


  sdffs1
  \DFF_1719/Q_reg 
  (
    .DIN(WX11654),
    .DIN_t(WX11654_t),
    .SDIN(CRC_OUT_1_22),
    .SDIN_t(CRC_OUT_1_22_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_23),
    .Q_t(CRC_OUT_1_23_t),
    .QN(n6301),
    .QN_t(n6301_t)
  );


  sdffs1
  \DFF_1718/Q_reg 
  (
    .DIN(WX11652),
    .DIN_t(WX11652_t),
    .SDIN(CRC_OUT_1_21),
    .SDIN_t(CRC_OUT_1_21_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_22),
    .Q_t(CRC_OUT_1_22_t),
    .QN(n6296),
    .QN_t(n6296_t)
  );


  sdffs1
  \DFF_1717/Q_reg 
  (
    .DIN(WX11650),
    .DIN_t(WX11650_t),
    .SDIN(CRC_OUT_1_20),
    .SDIN_t(CRC_OUT_1_20_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_21),
    .Q_t(CRC_OUT_1_21_t),
    .QN(n6291),
    .QN_t(n6291_t)
  );


  sdffs1
  \DFF_1716/Q_reg 
  (
    .DIN(WX11648),
    .DIN_t(WX11648_t),
    .SDIN(CRC_OUT_1_19),
    .SDIN_t(CRC_OUT_1_19_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_20),
    .Q_t(CRC_OUT_1_20_t),
    .QN(n6285),
    .QN_t(n6285_t)
  );


  sdffs1
  \DFF_1715/Q_reg 
  (
    .DIN(WX11646),
    .DIN_t(WX11646_t),
    .SDIN(CRC_OUT_1_18),
    .SDIN_t(CRC_OUT_1_18_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_19),
    .Q_t(CRC_OUT_1_19_t),
    .QN(n6280),
    .QN_t(n6280_t)
  );


  sdffs1
  \DFF_1714/Q_reg 
  (
    .DIN(WX11644),
    .DIN_t(WX11644_t),
    .SDIN(CRC_OUT_1_17),
    .SDIN_t(CRC_OUT_1_17_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_18),
    .Q_t(CRC_OUT_1_18_t),
    .QN(n6275),
    .QN_t(n6275_t)
  );


  sdffs1
  \DFF_1713/Q_reg 
  (
    .DIN(WX11642),
    .DIN_t(WX11642_t),
    .SDIN(CRC_OUT_1_16),
    .SDIN_t(CRC_OUT_1_16_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_17),
    .Q_t(CRC_OUT_1_17_t),
    .QN(n6270),
    .QN_t(n6270_t)
  );


  sdffs1
  \DFF_1712/Q_reg 
  (
    .DIN(WX11640),
    .DIN_t(WX11640_t),
    .SDIN(CRC_OUT_1_15),
    .SDIN_t(CRC_OUT_1_15_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_16),
    .Q_t(CRC_OUT_1_16_t),
    .QN(n6265),
    .QN_t(n6265_t)
  );


  sdffs1
  \DFF_1711/Q_reg 
  (
    .DIN(WX11638),
    .DIN_t(WX11638_t),
    .SDIN(CRC_OUT_1_14),
    .SDIN_t(CRC_OUT_1_14_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_15),
    .Q_t(CRC_OUT_1_15_t),
    .QN(n6260),
    .QN_t(n6260_t)
  );


  sdffs1
  \DFF_1710/Q_reg 
  (
    .DIN(WX11636),
    .DIN_t(WX11636_t),
    .SDIN(CRC_OUT_1_13),
    .SDIN_t(CRC_OUT_1_13_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_14),
    .Q_t(CRC_OUT_1_14_t),
    .QN(n6256),
    .QN_t(n6256_t)
  );


  sdffs1
  \DFF_1709/Q_reg 
  (
    .DIN(WX11634),
    .DIN_t(WX11634_t),
    .SDIN(CRC_OUT_1_12),
    .SDIN_t(CRC_OUT_1_12_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_13),
    .Q_t(CRC_OUT_1_13_t),
    .QN(n6252),
    .QN_t(n6252_t)
  );


  sdffs1
  \DFF_1708/Q_reg 
  (
    .DIN(WX11632),
    .DIN_t(WX11632_t),
    .SDIN(CRC_OUT_1_11),
    .SDIN_t(CRC_OUT_1_11_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_12),
    .Q_t(CRC_OUT_1_12_t),
    .QN(n6248),
    .QN_t(n6248_t)
  );


  sdffs1
  \DFF_1707/Q_reg 
  (
    .DIN(WX11630),
    .DIN_t(WX11630_t),
    .SDIN(CRC_OUT_1_10),
    .SDIN_t(CRC_OUT_1_10_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_11),
    .Q_t(CRC_OUT_1_11_t),
    .QN(n6244),
    .QN_t(n6244_t)
  );


  sdffs1
  \DFF_1706/Q_reg 
  (
    .DIN(WX11628),
    .DIN_t(WX11628_t),
    .SDIN(CRC_OUT_1_9),
    .SDIN_t(CRC_OUT_1_9_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_10),
    .Q_t(CRC_OUT_1_10_t),
    .QN(n6240),
    .QN_t(n6240_t)
  );


  sdffs1
  \DFF_1705/Q_reg 
  (
    .DIN(WX11626),
    .DIN_t(WX11626_t),
    .SDIN(CRC_OUT_1_8),
    .SDIN_t(CRC_OUT_1_8_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_9),
    .Q_t(CRC_OUT_1_9_t),
    .QN(n6236),
    .QN_t(n6236_t)
  );


  sdffs1
  \DFF_1704/Q_reg 
  (
    .DIN(WX11624),
    .DIN_t(WX11624_t),
    .SDIN(CRC_OUT_1_7),
    .SDIN_t(CRC_OUT_1_7_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_8),
    .Q_t(CRC_OUT_1_8_t),
    .QN(n6232),
    .QN_t(n6232_t)
  );


  sdffs1
  \DFF_1703/Q_reg 
  (
    .DIN(WX11622),
    .DIN_t(WX11622_t),
    .SDIN(CRC_OUT_1_6),
    .SDIN_t(CRC_OUT_1_6_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_7),
    .Q_t(CRC_OUT_1_7_t),
    .QN(n6228),
    .QN_t(n6228_t)
  );


  sdffs1
  \DFF_1702/Q_reg 
  (
    .DIN(WX11620),
    .DIN_t(WX11620_t),
    .SDIN(CRC_OUT_1_5),
    .SDIN_t(CRC_OUT_1_5_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_6),
    .Q_t(CRC_OUT_1_6_t),
    .QN(n6224),
    .QN_t(n6224_t)
  );


  sdffs1
  \DFF_1701/Q_reg 
  (
    .DIN(WX11618),
    .DIN_t(WX11618_t),
    .SDIN(CRC_OUT_1_4),
    .SDIN_t(CRC_OUT_1_4_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_5),
    .Q_t(CRC_OUT_1_5_t),
    .QN(n6220),
    .QN_t(n6220_t)
  );


  sdffs1
  \DFF_1700/Q_reg 
  (
    .DIN(WX11616),
    .DIN_t(WX11616_t),
    .SDIN(CRC_OUT_1_3),
    .SDIN_t(CRC_OUT_1_3_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_4),
    .Q_t(CRC_OUT_1_4_t),
    .QN(n6216),
    .QN_t(n6216_t)
  );


  sdffs1
  \DFF_1699/Q_reg 
  (
    .DIN(WX11614),
    .DIN_t(WX11614_t),
    .SDIN(CRC_OUT_1_2),
    .SDIN_t(CRC_OUT_1_2_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_3),
    .Q_t(CRC_OUT_1_3_t),
    .QN(n6212),
    .QN_t(n6212_t)
  );


  sdffs1
  \DFF_1698/Q_reg 
  (
    .DIN(WX11612),
    .DIN_t(WX11612_t),
    .SDIN(CRC_OUT_1_1),
    .SDIN_t(CRC_OUT_1_1_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_2),
    .Q_t(CRC_OUT_1_2_t),
    .QN(n6208),
    .QN_t(n6208_t)
  );


  sdffs1
  \DFF_1697/Q_reg 
  (
    .DIN(WX11610),
    .DIN_t(WX11610_t),
    .SDIN(CRC_OUT_1_0),
    .SDIN_t(CRC_OUT_1_0_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_1),
    .Q_t(CRC_OUT_1_1_t),
    .QN(n6204),
    .QN_t(n6204_t)
  );


  sdffs1
  \DFF_1696/Q_reg 
  (
    .DIN(WX11608),
    .DIN_t(WX11608_t),
    .SDIN(n7994),
    .SDIN_t(n7994_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_1_0),
    .Q_t(CRC_OUT_1_0_t),
    .QN(n6200),
    .QN_t(n6200_t)
  );


  sdffs1
  \DFF_1695/Q_reg 
  (
    .DIN(WX11242),
    .DIN_t(WX11242_t),
    .SDIN(n7993),
    .SDIN_t(n7993_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7994),
    .Q_t(n7994_t),
    .QN(n3317),
    .QN_t(n3317_t)
  );


  sdffs1
  \DFF_1694/Q_reg 
  (
    .DIN(WX11240),
    .DIN_t(WX11240_t),
    .SDIN(n7992),
    .SDIN_t(n7992_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7993),
    .Q_t(n7993_t),
    .QN(n3318),
    .QN_t(n3318_t)
  );


  sdffs1
  \DFF_1693/Q_reg 
  (
    .DIN(WX11238),
    .DIN_t(WX11238_t),
    .SDIN(n7991),
    .SDIN_t(n7991_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7992),
    .Q_t(n7992_t),
    .QN(n3319),
    .QN_t(n3319_t)
  );


  sdffs1
  \DFF_1692/Q_reg 
  (
    .DIN(WX11236),
    .DIN_t(WX11236_t),
    .SDIN(n7990),
    .SDIN_t(n7990_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7991),
    .Q_t(n7991_t),
    .QN(n3320),
    .QN_t(n3320_t)
  );


  sdffs1
  \DFF_1691/Q_reg 
  (
    .DIN(WX11234),
    .DIN_t(WX11234_t),
    .SDIN(n7989),
    .SDIN_t(n7989_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7990),
    .Q_t(n7990_t),
    .QN(n3321),
    .QN_t(n3321_t)
  );


  sdffs1
  \DFF_1690/Q_reg 
  (
    .DIN(WX11232),
    .DIN_t(WX11232_t),
    .SDIN(n7988),
    .SDIN_t(n7988_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7989),
    .Q_t(n7989_t),
    .QN(n3322),
    .QN_t(n3322_t)
  );


  sdffs1
  \DFF_1689/Q_reg 
  (
    .DIN(WX11230),
    .DIN_t(WX11230_t),
    .SDIN(n7987),
    .SDIN_t(n7987_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7988),
    .Q_t(n7988_t),
    .QN(n3323),
    .QN_t(n3323_t)
  );


  sdffs1
  \DFF_1688/Q_reg 
  (
    .DIN(WX11228),
    .DIN_t(WX11228_t),
    .SDIN(n7986),
    .SDIN_t(n7986_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7987),
    .Q_t(n7987_t),
    .QN(n3324),
    .QN_t(n3324_t)
  );


  sdffs1
  \DFF_1687/Q_reg 
  (
    .DIN(WX11226),
    .DIN_t(WX11226_t),
    .SDIN(n7985),
    .SDIN_t(n7985_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7986),
    .Q_t(n7986_t),
    .QN(n3325),
    .QN_t(n3325_t)
  );


  sdffs1
  \DFF_1686/Q_reg 
  (
    .DIN(WX11224),
    .DIN_t(WX11224_t),
    .SDIN(n7984),
    .SDIN_t(n7984_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7985),
    .Q_t(n7985_t),
    .QN(n3326),
    .QN_t(n3326_t)
  );


  sdffs1
  \DFF_1685/Q_reg 
  (
    .DIN(WX11222),
    .DIN_t(WX11222_t),
    .SDIN(n7983),
    .SDIN_t(n7983_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7984),
    .Q_t(n7984_t),
    .QN(n3327),
    .QN_t(n3327_t)
  );


  sdffs1
  \DFF_1684/Q_reg 
  (
    .DIN(WX11220),
    .DIN_t(WX11220_t),
    .SDIN(n7982),
    .SDIN_t(n7982_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7983),
    .Q_t(n7983_t),
    .QN(n3328),
    .QN_t(n3328_t)
  );


  sdffs1
  \DFF_1683/Q_reg 
  (
    .DIN(WX11218),
    .DIN_t(WX11218_t),
    .SDIN(n7981),
    .SDIN_t(n7981_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7982),
    .Q_t(n7982_t),
    .QN(n3329),
    .QN_t(n3329_t)
  );


  sdffs1
  \DFF_1682/Q_reg 
  (
    .DIN(WX11216),
    .DIN_t(WX11216_t),
    .SDIN(n7980),
    .SDIN_t(n7980_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7981),
    .Q_t(n7981_t),
    .QN(n3330),
    .QN_t(n3330_t)
  );


  sdffs1
  \DFF_1681/Q_reg 
  (
    .DIN(WX11214),
    .DIN_t(WX11214_t),
    .SDIN(n7979),
    .SDIN_t(n7979_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7980),
    .Q_t(n7980_t),
    .QN(n3331),
    .QN_t(n3331_t)
  );


  sdffs1
  \DFF_1680/Q_reg 
  (
    .DIN(WX11212),
    .DIN_t(WX11212_t),
    .SDIN(n7978),
    .SDIN_t(n7978_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7979),
    .Q_t(n7979_t),
    .QN(n3332),
    .QN_t(n3332_t)
  );


  sdffs1
  \DFF_1679/Q_reg 
  (
    .DIN(WX11210),
    .DIN_t(WX11210_t),
    .SDIN(n7977),
    .SDIN_t(n7977_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7978),
    .Q_t(n7978_t),
    .QN(n6264),
    .QN_t(n6264_t)
  );


  sdffs1
  \DFF_1678/Q_reg 
  (
    .DIN(WX11208),
    .DIN_t(WX11208_t),
    .SDIN(n7976),
    .SDIN_t(n7976_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7977),
    .Q_t(n7977_t),
    .QN(n6269),
    .QN_t(n6269_t)
  );


  sdffs1
  \DFF_1677/Q_reg 
  (
    .DIN(WX11206),
    .DIN_t(WX11206_t),
    .SDIN(n7975),
    .SDIN_t(n7975_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7976),
    .Q_t(n7976_t),
    .QN(n6274),
    .QN_t(n6274_t)
  );


  sdffs1
  \DFF_1676/Q_reg 
  (
    .DIN(WX11204),
    .DIN_t(WX11204_t),
    .SDIN(n7974),
    .SDIN_t(n7974_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7975),
    .Q_t(n7975_t),
    .QN(n6279),
    .QN_t(n6279_t)
  );


  sdffs1
  \DFF_1675/Q_reg 
  (
    .DIN(WX11202),
    .DIN_t(WX11202_t),
    .SDIN(n7973),
    .SDIN_t(n7973_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7974),
    .Q_t(n7974_t),
    .QN(n6284),
    .QN_t(n6284_t)
  );


  sdffs1
  \DFF_1674/Q_reg 
  (
    .DIN(WX11200),
    .DIN_t(WX11200_t),
    .SDIN(n7972),
    .SDIN_t(n7972_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7973),
    .Q_t(n7973_t),
    .QN(n6290),
    .QN_t(n6290_t)
  );


  sdffs1
  \DFF_1673/Q_reg 
  (
    .DIN(WX11198),
    .DIN_t(WX11198_t),
    .SDIN(n7971),
    .SDIN_t(n7971_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7972),
    .Q_t(n7972_t),
    .QN(n6295),
    .QN_t(n6295_t)
  );


  sdffs1
  \DFF_1672/Q_reg 
  (
    .DIN(WX11196),
    .DIN_t(WX11196_t),
    .SDIN(n7970),
    .SDIN_t(n7970_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7971),
    .Q_t(n7971_t),
    .QN(n6300),
    .QN_t(n6300_t)
  );


  sdffs1
  \DFF_1671/Q_reg 
  (
    .DIN(WX11194),
    .DIN_t(WX11194_t),
    .SDIN(n7969),
    .SDIN_t(n7969_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7970),
    .Q_t(n7970_t),
    .QN(n6305),
    .QN_t(n6305_t)
  );


  sdffs1
  \DFF_1670/Q_reg 
  (
    .DIN(WX11192),
    .DIN_t(WX11192_t),
    .SDIN(n7968),
    .SDIN_t(n7968_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7969),
    .Q_t(n7969_t),
    .QN(n6310),
    .QN_t(n6310_t)
  );


  sdffs1
  \DFF_1669/Q_reg 
  (
    .DIN(WX11190),
    .DIN_t(WX11190_t),
    .SDIN(n7967),
    .SDIN_t(n7967_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7968),
    .Q_t(n7968_t),
    .QN(n6315),
    .QN_t(n6315_t)
  );


  sdffs1
  \DFF_1668/Q_reg 
  (
    .DIN(WX11188),
    .DIN_t(WX11188_t),
    .SDIN(n7966),
    .SDIN_t(n7966_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7967),
    .Q_t(n7967_t),
    .QN(n6320),
    .QN_t(n6320_t)
  );


  sdffs1
  \DFF_1667/Q_reg 
  (
    .DIN(WX11186),
    .DIN_t(WX11186_t),
    .SDIN(n7965),
    .SDIN_t(n7965_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7966),
    .Q_t(n7966_t),
    .QN(n6325),
    .QN_t(n6325_t)
  );


  sdffs1
  \DFF_1666/Q_reg 
  (
    .DIN(WX11184),
    .DIN_t(WX11184_t),
    .SDIN(n7964),
    .SDIN_t(n7964_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7965),
    .Q_t(n7965_t),
    .QN(n6330),
    .QN_t(n6330_t)
  );


  sdffs1
  \DFF_1665/Q_reg 
  (
    .DIN(WX11182),
    .DIN_t(WX11182_t),
    .SDIN(n7963),
    .SDIN_t(n7963_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7964),
    .Q_t(n7964_t),
    .QN(n6335),
    .QN_t(n6335_t)
  );


  sdffs1
  \DFF_1664/Q_reg 
  (
    .DIN(WX11180),
    .DIN_t(WX11180_t),
    .SDIN(n7962),
    .SDIN_t(n7962_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7963),
    .Q_t(n7963_t),
    .QN(n6341),
    .QN_t(n6341_t)
  );


  sdffs1
  \DFF_1663/Q_reg 
  (
    .DIN(WX11178),
    .DIN_t(WX11178_t),
    .SDIN(n7961),
    .SDIN_t(n7961_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7962),
    .Q_t(n7962_t),
    .QN(n6199),
    .QN_t(n6199_t)
  );


  sdffs1
  \DFF_1662/Q_reg 
  (
    .DIN(WX11176),
    .DIN_t(WX11176_t),
    .SDIN(n7960),
    .SDIN_t(n7960_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7961),
    .Q_t(n7961_t),
    .QN(n6203),
    .QN_t(n6203_t)
  );


  sdffs1
  \DFF_1661/Q_reg 
  (
    .DIN(WX11174),
    .DIN_t(WX11174_t),
    .SDIN(n7959),
    .SDIN_t(n7959_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7960),
    .Q_t(n7960_t),
    .QN(n6207),
    .QN_t(n6207_t)
  );


  sdffs1
  \DFF_1660/Q_reg 
  (
    .DIN(WX11172),
    .DIN_t(WX11172_t),
    .SDIN(n7958),
    .SDIN_t(n7958_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7959),
    .Q_t(n7959_t),
    .QN(n6211),
    .QN_t(n6211_t)
  );


  sdffs1
  \DFF_1659/Q_reg 
  (
    .DIN(WX11170),
    .DIN_t(WX11170_t),
    .SDIN(n7957),
    .SDIN_t(n7957_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7958),
    .Q_t(n7958_t),
    .QN(n6215),
    .QN_t(n6215_t)
  );


  sdffs1
  \DFF_1658/Q_reg 
  (
    .DIN(WX11168),
    .DIN_t(WX11168_t),
    .SDIN(n7956),
    .SDIN_t(n7956_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7957),
    .Q_t(n7957_t),
    .QN(n6219),
    .QN_t(n6219_t)
  );


  sdffs1
  \DFF_1657/Q_reg 
  (
    .DIN(WX11166),
    .DIN_t(WX11166_t),
    .SDIN(n7955),
    .SDIN_t(n7955_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7956),
    .Q_t(n7956_t),
    .QN(n6223),
    .QN_t(n6223_t)
  );


  sdffs1
  \DFF_1656/Q_reg 
  (
    .DIN(WX11164),
    .DIN_t(WX11164_t),
    .SDIN(n7954),
    .SDIN_t(n7954_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7955),
    .Q_t(n7955_t),
    .QN(n6227),
    .QN_t(n6227_t)
  );


  sdffs1
  \DFF_1655/Q_reg 
  (
    .DIN(WX11162),
    .DIN_t(WX11162_t),
    .SDIN(n7953),
    .SDIN_t(n7953_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7954),
    .Q_t(n7954_t),
    .QN(n6231),
    .QN_t(n6231_t)
  );


  sdffs1
  \DFF_1654/Q_reg 
  (
    .DIN(WX11160),
    .DIN_t(WX11160_t),
    .SDIN(n7952),
    .SDIN_t(n7952_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7953),
    .Q_t(n7953_t),
    .QN(n6235),
    .QN_t(n6235_t)
  );


  sdffs1
  \DFF_1653/Q_reg 
  (
    .DIN(WX11158),
    .DIN_t(WX11158_t),
    .SDIN(n7951),
    .SDIN_t(n7951_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7952),
    .Q_t(n7952_t),
    .QN(n6239),
    .QN_t(n6239_t)
  );


  sdffs1
  \DFF_1652/Q_reg 
  (
    .DIN(WX11156),
    .DIN_t(WX11156_t),
    .SDIN(n7950),
    .SDIN_t(n7950_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7951),
    .Q_t(n7951_t),
    .QN(n6243),
    .QN_t(n6243_t)
  );


  sdffs1
  \DFF_1651/Q_reg 
  (
    .DIN(WX11154),
    .DIN_t(WX11154_t),
    .SDIN(n7949),
    .SDIN_t(n7949_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7950),
    .Q_t(n7950_t),
    .QN(n6247),
    .QN_t(n6247_t)
  );


  sdffs1
  \DFF_1650/Q_reg 
  (
    .DIN(WX11152),
    .DIN_t(WX11152_t),
    .SDIN(n7948),
    .SDIN_t(n7948_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7949),
    .Q_t(n7949_t),
    .QN(n6251),
    .QN_t(n6251_t)
  );


  sdffs1
  \DFF_1649/Q_reg 
  (
    .DIN(WX11150),
    .DIN_t(WX11150_t),
    .SDIN(n7947),
    .SDIN_t(n7947_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7948),
    .Q_t(n7948_t),
    .QN(n6255),
    .QN_t(n6255_t)
  );


  sdffs1
  \DFF_1648/Q_reg 
  (
    .DIN(WX11148),
    .DIN_t(WX11148_t),
    .SDIN(n7946),
    .SDIN_t(n7946_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7947),
    .Q_t(n7947_t),
    .QN(n6259),
    .QN_t(n6259_t)
  );


  sdffs1
  \DFF_1647/Q_reg 
  (
    .DIN(WX11146),
    .DIN_t(WX11146_t),
    .SDIN(n7945),
    .SDIN_t(n7945_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7946),
    .Q_t(n7946_t),
    .QN(n6263),
    .QN_t(n6263_t)
  );


  sdffs1
  \DFF_1646/Q_reg 
  (
    .DIN(WX11144),
    .DIN_t(WX11144_t),
    .SDIN(n7944),
    .SDIN_t(n7944_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7945),
    .Q_t(n7945_t),
    .QN(n6268),
    .QN_t(n6268_t)
  );


  sdffs1
  \DFF_1645/Q_reg 
  (
    .DIN(WX11142),
    .DIN_t(WX11142_t),
    .SDIN(n7943),
    .SDIN_t(n7943_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7944),
    .Q_t(n7944_t),
    .QN(n6273),
    .QN_t(n6273_t)
  );


  sdffs1
  \DFF_1644/Q_reg 
  (
    .DIN(WX11140),
    .DIN_t(WX11140_t),
    .SDIN(n7942),
    .SDIN_t(n7942_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7943),
    .Q_t(n7943_t),
    .QN(n6278),
    .QN_t(n6278_t)
  );


  sdffs1
  \DFF_1643/Q_reg 
  (
    .DIN(WX11138),
    .DIN_t(WX11138_t),
    .SDIN(n7941),
    .SDIN_t(n7941_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7942),
    .Q_t(n7942_t),
    .QN(n6283),
    .QN_t(n6283_t)
  );


  sdffs1
  \DFF_1642/Q_reg 
  (
    .DIN(WX11136),
    .DIN_t(WX11136_t),
    .SDIN(n7940),
    .SDIN_t(n7940_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7941),
    .Q_t(n7941_t),
    .QN(n6289),
    .QN_t(n6289_t)
  );


  sdffs1
  \DFF_1641/Q_reg 
  (
    .DIN(WX11134),
    .DIN_t(WX11134_t),
    .SDIN(n7939),
    .SDIN_t(n7939_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7940),
    .Q_t(n7940_t),
    .QN(n6294),
    .QN_t(n6294_t)
  );


  sdffs1
  \DFF_1640/Q_reg 
  (
    .DIN(WX11132),
    .DIN_t(WX11132_t),
    .SDIN(n7938),
    .SDIN_t(n7938_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7939),
    .Q_t(n7939_t),
    .QN(n6299),
    .QN_t(n6299_t)
  );


  sdffs1
  \DFF_1639/Q_reg 
  (
    .DIN(WX11130),
    .DIN_t(WX11130_t),
    .SDIN(n7937),
    .SDIN_t(n7937_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7938),
    .Q_t(n7938_t),
    .QN(n6304),
    .QN_t(n6304_t)
  );


  sdffs1
  \DFF_1638/Q_reg 
  (
    .DIN(WX11128),
    .DIN_t(WX11128_t),
    .SDIN(n7936),
    .SDIN_t(n7936_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7937),
    .Q_t(n7937_t),
    .QN(n6309),
    .QN_t(n6309_t)
  );


  sdffs1
  \DFF_1637/Q_reg 
  (
    .DIN(WX11126),
    .DIN_t(WX11126_t),
    .SDIN(n7935),
    .SDIN_t(n7935_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7936),
    .Q_t(n7936_t),
    .QN(n6314),
    .QN_t(n6314_t)
  );


  sdffs1
  \DFF_1636/Q_reg 
  (
    .DIN(WX11124),
    .DIN_t(WX11124_t),
    .SDIN(n7934),
    .SDIN_t(n7934_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7935),
    .Q_t(n7935_t),
    .QN(n6319),
    .QN_t(n6319_t)
  );


  sdffs1
  \DFF_1635/Q_reg 
  (
    .DIN(WX11122),
    .DIN_t(WX11122_t),
    .SDIN(n7933),
    .SDIN_t(n7933_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7934),
    .Q_t(n7934_t),
    .QN(n6324),
    .QN_t(n6324_t)
  );


  sdffs1
  \DFF_1634/Q_reg 
  (
    .DIN(WX11120),
    .DIN_t(WX11120_t),
    .SDIN(n7932),
    .SDIN_t(n7932_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7933),
    .Q_t(n7933_t),
    .QN(n6329),
    .QN_t(n6329_t)
  );


  sdffs1
  \DFF_1633/Q_reg 
  (
    .DIN(WX11118),
    .DIN_t(WX11118_t),
    .SDIN(n7931),
    .SDIN_t(n7931_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7932),
    .Q_t(n7932_t),
    .QN(n6334),
    .QN_t(n6334_t)
  );


  sdffs1
  \DFF_1632/Q_reg 
  (
    .DIN(WX11116),
    .DIN_t(WX11116_t),
    .SDIN(n6198),
    .SDIN_t(n6198_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7931),
    .Q_t(n7931_t),
    .QN(n6340),
    .QN_t(n6340_t)
  );


  sdffs1
  \DFF_1631/Q_reg 
  (
    .DIN(WX11114),
    .DIN_t(WX11114_t),
    .SDIN(n6202),
    .SDIN_t(n6202_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6198),
    .Q_t(n6198_t)
  );


  sdffs1
  \DFF_1630/Q_reg 
  (
    .DIN(WX11112),
    .DIN_t(WX11112_t),
    .SDIN(n6206),
    .SDIN_t(n6206_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6202),
    .Q_t(n6202_t)
  );


  sdffs1
  \DFF_1629/Q_reg 
  (
    .DIN(WX11110),
    .DIN_t(WX11110_t),
    .SDIN(n6210),
    .SDIN_t(n6210_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6206),
    .Q_t(n6206_t)
  );


  sdffs1
  \DFF_1628/Q_reg 
  (
    .DIN(WX11108),
    .DIN_t(WX11108_t),
    .SDIN(n6214),
    .SDIN_t(n6214_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6210),
    .Q_t(n6210_t)
  );


  sdffs1
  \DFF_1627/Q_reg 
  (
    .DIN(WX11106),
    .DIN_t(WX11106_t),
    .SDIN(n6218),
    .SDIN_t(n6218_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6214),
    .Q_t(n6214_t)
  );


  sdffs1
  \DFF_1626/Q_reg 
  (
    .DIN(WX11104),
    .DIN_t(WX11104_t),
    .SDIN(n6222),
    .SDIN_t(n6222_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6218),
    .Q_t(n6218_t)
  );


  sdffs1
  \DFF_1625/Q_reg 
  (
    .DIN(WX11102),
    .DIN_t(WX11102_t),
    .SDIN(n6226),
    .SDIN_t(n6226_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6222),
    .Q_t(n6222_t)
  );


  sdffs1
  \DFF_1624/Q_reg 
  (
    .DIN(WX11100),
    .DIN_t(WX11100_t),
    .SDIN(n6230),
    .SDIN_t(n6230_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6226),
    .Q_t(n6226_t)
  );


  sdffs1
  \DFF_1623/Q_reg 
  (
    .DIN(WX11098),
    .DIN_t(WX11098_t),
    .SDIN(n6234),
    .SDIN_t(n6234_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6230),
    .Q_t(n6230_t)
  );


  sdffs1
  \DFF_1622/Q_reg 
  (
    .DIN(WX11096),
    .DIN_t(WX11096_t),
    .SDIN(n6238),
    .SDIN_t(n6238_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6234),
    .Q_t(n6234_t)
  );


  sdffs1
  \DFF_1621/Q_reg 
  (
    .DIN(WX11094),
    .DIN_t(WX11094_t),
    .SDIN(n6242),
    .SDIN_t(n6242_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6238),
    .Q_t(n6238_t)
  );


  sdffs1
  \DFF_1620/Q_reg 
  (
    .DIN(WX11092),
    .DIN_t(WX11092_t),
    .SDIN(n6246),
    .SDIN_t(n6246_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6242),
    .Q_t(n6242_t)
  );


  sdffs1
  \DFF_1619/Q_reg 
  (
    .DIN(WX11090),
    .DIN_t(WX11090_t),
    .SDIN(n6250),
    .SDIN_t(n6250_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6246),
    .Q_t(n6246_t)
  );


  sdffs1
  \DFF_1618/Q_reg 
  (
    .DIN(WX11088),
    .DIN_t(WX11088_t),
    .SDIN(n6254),
    .SDIN_t(n6254_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6250),
    .Q_t(n6250_t)
  );


  sdffs1
  \DFF_1617/Q_reg 
  (
    .DIN(WX11086),
    .DIN_t(WX11086_t),
    .SDIN(n6258),
    .SDIN_t(n6258_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6254),
    .Q_t(n6254_t)
  );


  sdffs1
  \DFF_1616/Q_reg 
  (
    .DIN(WX11084),
    .DIN_t(WX11084_t),
    .SDIN(n6262),
    .SDIN_t(n6262_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6258),
    .Q_t(n6258_t)
  );


  sdffs1
  \DFF_1615/Q_reg 
  (
    .DIN(WX11082),
    .DIN_t(WX11082_t),
    .SDIN(n6267),
    .SDIN_t(n6267_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6262),
    .Q_t(n6262_t)
  );


  sdffs1
  \DFF_1614/Q_reg 
  (
    .DIN(WX11080),
    .DIN_t(WX11080_t),
    .SDIN(n6272),
    .SDIN_t(n6272_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6267),
    .Q_t(n6267_t)
  );


  sdffs1
  \DFF_1613/Q_reg 
  (
    .DIN(WX11078),
    .DIN_t(WX11078_t),
    .SDIN(n6277),
    .SDIN_t(n6277_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6272),
    .Q_t(n6272_t)
  );


  sdffs1
  \DFF_1612/Q_reg 
  (
    .DIN(WX11076),
    .DIN_t(WX11076_t),
    .SDIN(n6282),
    .SDIN_t(n6282_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6277),
    .Q_t(n6277_t)
  );


  sdffs1
  \DFF_1611/Q_reg 
  (
    .DIN(WX11074),
    .DIN_t(WX11074_t),
    .SDIN(n6288),
    .SDIN_t(n6288_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6282),
    .Q_t(n6282_t)
  );


  sdffs1
  \DFF_1610/Q_reg 
  (
    .DIN(WX11072),
    .DIN_t(WX11072_t),
    .SDIN(n6293),
    .SDIN_t(n6293_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6288),
    .Q_t(n6288_t)
  );


  sdffs1
  \DFF_1609/Q_reg 
  (
    .DIN(WX11070),
    .DIN_t(WX11070_t),
    .SDIN(n6298),
    .SDIN_t(n6298_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6293),
    .Q_t(n6293_t)
  );


  sdffs1
  \DFF_1608/Q_reg 
  (
    .DIN(WX11068),
    .DIN_t(WX11068_t),
    .SDIN(n6303),
    .SDIN_t(n6303_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6298),
    .Q_t(n6298_t)
  );


  sdffs1
  \DFF_1607/Q_reg 
  (
    .DIN(WX11066),
    .DIN_t(WX11066_t),
    .SDIN(n6308),
    .SDIN_t(n6308_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6303),
    .Q_t(n6303_t)
  );


  sdffs1
  \DFF_1606/Q_reg 
  (
    .DIN(WX11064),
    .DIN_t(WX11064_t),
    .SDIN(n6313),
    .SDIN_t(n6313_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6308),
    .Q_t(n6308_t)
  );


  sdffs1
  \DFF_1605/Q_reg 
  (
    .DIN(WX11062),
    .DIN_t(WX11062_t),
    .SDIN(n6318),
    .SDIN_t(n6318_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6313),
    .Q_t(n6313_t)
  );


  sdffs1
  \DFF_1604/Q_reg 
  (
    .DIN(WX11060),
    .DIN_t(WX11060_t),
    .SDIN(n6323),
    .SDIN_t(n6323_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6318),
    .Q_t(n6318_t)
  );


  sdffs1
  \DFF_1603/Q_reg 
  (
    .DIN(WX11058),
    .DIN_t(WX11058_t),
    .SDIN(n6328),
    .SDIN_t(n6328_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6323),
    .Q_t(n6323_t)
  );


  sdffs1
  \DFF_1602/Q_reg 
  (
    .DIN(WX11056),
    .DIN_t(WX11056_t),
    .SDIN(n6333),
    .SDIN_t(n6333_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6328),
    .Q_t(n6328_t)
  );


  sdffs1
  \DFF_1601/Q_reg 
  (
    .DIN(WX11054),
    .DIN_t(WX11054_t),
    .SDIN(n6339),
    .SDIN_t(n6339_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6333),
    .Q_t(n6333_t)
  );


  sdffs1
  \DFF_1600/Q_reg 
  (
    .DIN(WX11052),
    .DIN_t(WX11052_t),
    .SDIN(n7930),
    .SDIN_t(n7930_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6339),
    .Q_t(n6339_t)
  );


  sdffs1
  \DFF_1599/Q_reg 
  (
    .DIN(WX11050),
    .DIN_t(WX11050_t),
    .SDIN(n7929),
    .SDIN_t(n7929_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7930),
    .Q_t(n7930_t),
    .QN(n6197),
    .QN_t(n6197_t)
  );


  sdffs1
  \DFF_1598/Q_reg 
  (
    .DIN(WX11048),
    .DIN_t(WX11048_t),
    .SDIN(n7928),
    .SDIN_t(n7928_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7929),
    .Q_t(n7929_t),
    .QN(n6201),
    .QN_t(n6201_t)
  );


  sdffs1
  \DFF_1597/Q_reg 
  (
    .DIN(WX11046),
    .DIN_t(WX11046_t),
    .SDIN(n7927),
    .SDIN_t(n7927_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7928),
    .Q_t(n7928_t),
    .QN(n6205),
    .QN_t(n6205_t)
  );


  sdffs1
  \DFF_1596/Q_reg 
  (
    .DIN(WX11044),
    .DIN_t(WX11044_t),
    .SDIN(n7926),
    .SDIN_t(n7926_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7927),
    .Q_t(n7927_t),
    .QN(n6209),
    .QN_t(n6209_t)
  );


  sdffs1
  \DFF_1595/Q_reg 
  (
    .DIN(WX11042),
    .DIN_t(WX11042_t),
    .SDIN(n7925),
    .SDIN_t(n7925_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7926),
    .Q_t(n7926_t),
    .QN(n6213),
    .QN_t(n6213_t)
  );


  sdffs1
  \DFF_1594/Q_reg 
  (
    .DIN(WX11040),
    .DIN_t(WX11040_t),
    .SDIN(n7924),
    .SDIN_t(n7924_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7925),
    .Q_t(n7925_t),
    .QN(n6217),
    .QN_t(n6217_t)
  );


  sdffs1
  \DFF_1593/Q_reg 
  (
    .DIN(WX11038),
    .DIN_t(WX11038_t),
    .SDIN(n7923),
    .SDIN_t(n7923_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7924),
    .Q_t(n7924_t),
    .QN(n6221),
    .QN_t(n6221_t)
  );


  sdffs1
  \DFF_1592/Q_reg 
  (
    .DIN(WX11036),
    .DIN_t(WX11036_t),
    .SDIN(n7922),
    .SDIN_t(n7922_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7923),
    .Q_t(n7923_t),
    .QN(n6225),
    .QN_t(n6225_t)
  );


  sdffs1
  \DFF_1591/Q_reg 
  (
    .DIN(WX11034),
    .DIN_t(WX11034_t),
    .SDIN(n7921),
    .SDIN_t(n7921_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7922),
    .Q_t(n7922_t),
    .QN(n6229),
    .QN_t(n6229_t)
  );


  sdffs1
  \DFF_1590/Q_reg 
  (
    .DIN(WX11032),
    .DIN_t(WX11032_t),
    .SDIN(n7920),
    .SDIN_t(n7920_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7921),
    .Q_t(n7921_t),
    .QN(n6233),
    .QN_t(n6233_t)
  );


  sdffs1
  \DFF_1589/Q_reg 
  (
    .DIN(WX11030),
    .DIN_t(WX11030_t),
    .SDIN(n7919),
    .SDIN_t(n7919_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7920),
    .Q_t(n7920_t),
    .QN(n6237),
    .QN_t(n6237_t)
  );


  sdffs1
  \DFF_1588/Q_reg 
  (
    .DIN(WX11028),
    .DIN_t(WX11028_t),
    .SDIN(n7918),
    .SDIN_t(n7918_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7919),
    .Q_t(n7919_t),
    .QN(n6241),
    .QN_t(n6241_t)
  );


  sdffs1
  \DFF_1587/Q_reg 
  (
    .DIN(WX11026),
    .DIN_t(WX11026_t),
    .SDIN(n7917),
    .SDIN_t(n7917_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7918),
    .Q_t(n7918_t),
    .QN(n6245),
    .QN_t(n6245_t)
  );


  sdffs1
  \DFF_1586/Q_reg 
  (
    .DIN(WX11024),
    .DIN_t(WX11024_t),
    .SDIN(n7916),
    .SDIN_t(n7916_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7917),
    .Q_t(n7917_t),
    .QN(n6249),
    .QN_t(n6249_t)
  );


  sdffs1
  \DFF_1585/Q_reg 
  (
    .DIN(WX11022),
    .DIN_t(WX11022_t),
    .SDIN(n7915),
    .SDIN_t(n7915_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7916),
    .Q_t(n7916_t),
    .QN(n6253),
    .QN_t(n6253_t)
  );


  sdffs1
  \DFF_1584/Q_reg 
  (
    .DIN(WX11020),
    .DIN_t(WX11020_t),
    .SDIN(n7914),
    .SDIN_t(n7914_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7915),
    .Q_t(n7915_t),
    .QN(n6257),
    .QN_t(n6257_t)
  );


  sdffs1
  \DFF_1583/Q_reg 
  (
    .DIN(WX11018),
    .DIN_t(WX11018_t),
    .SDIN(n7913),
    .SDIN_t(n7913_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7914),
    .Q_t(n7914_t),
    .QN(n6261),
    .QN_t(n6261_t)
  );


  sdffs1
  \DFF_1582/Q_reg 
  (
    .DIN(WX11016),
    .DIN_t(WX11016_t),
    .SDIN(n7912),
    .SDIN_t(n7912_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7913),
    .Q_t(n7913_t),
    .QN(n6266),
    .QN_t(n6266_t)
  );


  sdffs1
  \DFF_1581/Q_reg 
  (
    .DIN(WX11014),
    .DIN_t(WX11014_t),
    .SDIN(n7911),
    .SDIN_t(n7911_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7912),
    .Q_t(n7912_t),
    .QN(n6271),
    .QN_t(n6271_t)
  );


  sdffs1
  \DFF_1580/Q_reg 
  (
    .DIN(WX11012),
    .DIN_t(WX11012_t),
    .SDIN(n7910),
    .SDIN_t(n7910_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7911),
    .Q_t(n7911_t),
    .QN(n6276),
    .QN_t(n6276_t)
  );


  sdffs1
  \DFF_1579/Q_reg 
  (
    .DIN(WX11010),
    .DIN_t(WX11010_t),
    .SDIN(n7909),
    .SDIN_t(n7909_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7910),
    .Q_t(n7910_t),
    .QN(n6281),
    .QN_t(n6281_t)
  );


  sdffs1
  \DFF_1578/Q_reg 
  (
    .DIN(WX11008),
    .DIN_t(WX11008_t),
    .SDIN(n7908),
    .SDIN_t(n7908_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7909),
    .Q_t(n7909_t),
    .QN(n6287),
    .QN_t(n6287_t)
  );


  sdffs1
  \DFF_1577/Q_reg 
  (
    .DIN(WX11006),
    .DIN_t(WX11006_t),
    .SDIN(n7907),
    .SDIN_t(n7907_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7908),
    .Q_t(n7908_t),
    .QN(n6292),
    .QN_t(n6292_t)
  );


  sdffs1
  \DFF_1576/Q_reg 
  (
    .DIN(WX11004),
    .DIN_t(WX11004_t),
    .SDIN(n7906),
    .SDIN_t(n7906_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7907),
    .Q_t(n7907_t),
    .QN(n6297),
    .QN_t(n6297_t)
  );


  sdffs1
  \DFF_1575/Q_reg 
  (
    .DIN(WX11002),
    .DIN_t(WX11002_t),
    .SDIN(n7905),
    .SDIN_t(n7905_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7906),
    .Q_t(n7906_t),
    .QN(n6302),
    .QN_t(n6302_t)
  );


  sdffs1
  \DFF_1574/Q_reg 
  (
    .DIN(WX11000),
    .DIN_t(WX11000_t),
    .SDIN(n7904),
    .SDIN_t(n7904_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7905),
    .Q_t(n7905_t),
    .QN(n6307),
    .QN_t(n6307_t)
  );


  sdffs1
  \DFF_1573/Q_reg 
  (
    .DIN(WX10998),
    .DIN_t(WX10998_t),
    .SDIN(n7903),
    .SDIN_t(n7903_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7904),
    .Q_t(n7904_t),
    .QN(n6312),
    .QN_t(n6312_t)
  );


  sdffs1
  \DFF_1572/Q_reg 
  (
    .DIN(WX10996),
    .DIN_t(WX10996_t),
    .SDIN(n7902),
    .SDIN_t(n7902_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7903),
    .Q_t(n7903_t),
    .QN(n6317),
    .QN_t(n6317_t)
  );


  sdffs1
  \DFF_1571/Q_reg 
  (
    .DIN(WX10994),
    .DIN_t(WX10994_t),
    .SDIN(n7901),
    .SDIN_t(n7901_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7902),
    .Q_t(n7902_t),
    .QN(n6322),
    .QN_t(n6322_t)
  );


  sdffs1
  \DFF_1570/Q_reg 
  (
    .DIN(WX10992),
    .DIN_t(WX10992_t),
    .SDIN(n7900),
    .SDIN_t(n7900_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7901),
    .Q_t(n7901_t),
    .QN(n6327),
    .QN_t(n6327_t)
  );


  sdffs1
  \DFF_1569/Q_reg 
  (
    .DIN(WX10990),
    .DIN_t(WX10990_t),
    .SDIN(n7899),
    .SDIN_t(n7899_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7900),
    .Q_t(n7900_t),
    .QN(n6332),
    .QN_t(n6332_t)
  );


  sdffs1
  \DFF_1568/Q_reg 
  (
    .DIN(WX10988),
    .DIN_t(WX10988_t),
    .SDIN(n7898),
    .SDIN_t(n7898_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7899),
    .Q_t(n7899_t),
    .QN(n6338),
    .QN_t(n6338_t)
  );


  sdffs1
  \DFF_1567/Q_reg 
  (
    .DIN(WX10890),
    .DIN_t(WX10890_t),
    .SDIN(n7897),
    .SDIN_t(n7897_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7898),
    .Q_t(n7898_t),
    .QN(n6344),
    .QN_t(n6344_t)
  );


  sdffs1
  \DFF_1566/Q_reg 
  (
    .DIN(WX10888),
    .DIN_t(WX10888_t),
    .SDIN(n7896),
    .SDIN_t(n7896_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7897),
    .Q_t(n7897_t),
    .QN(n6345),
    .QN_t(n6345_t)
  );


  sdffs1
  \DFF_1565/Q_reg 
  (
    .DIN(WX10886),
    .DIN_t(WX10886_t),
    .SDIN(n7895),
    .SDIN_t(n7895_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7896),
    .Q_t(n7896_t),
    .QN(n6346),
    .QN_t(n6346_t)
  );


  sdffs1
  \DFF_1564/Q_reg 
  (
    .DIN(WX10884),
    .DIN_t(WX10884_t),
    .SDIN(n7894),
    .SDIN_t(n7894_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7895),
    .Q_t(n7895_t),
    .QN(n6347),
    .QN_t(n6347_t)
  );


  sdffs1
  \DFF_1563/Q_reg 
  (
    .DIN(WX10882),
    .DIN_t(WX10882_t),
    .SDIN(n7893),
    .SDIN_t(n7893_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7894),
    .Q_t(n7894_t),
    .QN(n6348),
    .QN_t(n6348_t)
  );


  sdffs1
  \DFF_1562/Q_reg 
  (
    .DIN(WX10880),
    .DIN_t(WX10880_t),
    .SDIN(n7892),
    .SDIN_t(n7892_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7893),
    .Q_t(n7893_t),
    .QN(n6349),
    .QN_t(n6349_t)
  );


  sdffs1
  \DFF_1561/Q_reg 
  (
    .DIN(WX10878),
    .DIN_t(WX10878_t),
    .SDIN(n7891),
    .SDIN_t(n7891_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7892),
    .Q_t(n7892_t),
    .QN(n6350),
    .QN_t(n6350_t)
  );


  sdffs1
  \DFF_1560/Q_reg 
  (
    .DIN(WX10876),
    .DIN_t(WX10876_t),
    .SDIN(n7890),
    .SDIN_t(n7890_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7891),
    .Q_t(n7891_t),
    .QN(n6351),
    .QN_t(n6351_t)
  );


  sdffs1
  \DFF_1559/Q_reg 
  (
    .DIN(WX10874),
    .DIN_t(WX10874_t),
    .SDIN(n7889),
    .SDIN_t(n7889_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7890),
    .Q_t(n7890_t),
    .QN(n6352),
    .QN_t(n6352_t)
  );


  sdffs1
  \DFF_1558/Q_reg 
  (
    .DIN(WX10872),
    .DIN_t(WX10872_t),
    .SDIN(n7888),
    .SDIN_t(n7888_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7889),
    .Q_t(n7889_t),
    .QN(n6353),
    .QN_t(n6353_t)
  );


  sdffs1
  \DFF_1557/Q_reg 
  (
    .DIN(WX10870),
    .DIN_t(WX10870_t),
    .SDIN(n7887),
    .SDIN_t(n7887_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7888),
    .Q_t(n7888_t),
    .QN(n6355),
    .QN_t(n6355_t)
  );


  sdffs1
  \DFF_1556/Q_reg 
  (
    .DIN(WX10868),
    .DIN_t(WX10868_t),
    .SDIN(n7886),
    .SDIN_t(n7886_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7887),
    .Q_t(n7887_t),
    .QN(n6356),
    .QN_t(n6356_t)
  );


  sdffs1
  \DFF_1555/Q_reg 
  (
    .DIN(WX10866),
    .DIN_t(WX10866_t),
    .SDIN(n7885),
    .SDIN_t(n7885_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7886),
    .Q_t(n7886_t),
    .QN(n6357),
    .QN_t(n6357_t)
  );


  sdffs1
  \DFF_1554/Q_reg 
  (
    .DIN(WX10864),
    .DIN_t(WX10864_t),
    .SDIN(n7884),
    .SDIN_t(n7884_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7885),
    .Q_t(n7885_t),
    .QN(n6358),
    .QN_t(n6358_t)
  );


  sdffs1
  \DFF_1553/Q_reg 
  (
    .DIN(WX10862),
    .DIN_t(WX10862_t),
    .SDIN(n7883),
    .SDIN_t(n7883_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7884),
    .Q_t(n7884_t),
    .QN(n6359),
    .QN_t(n6359_t)
  );


  sdffs1
  \DFF_1552/Q_reg 
  (
    .DIN(WX10860),
    .DIN_t(WX10860_t),
    .SDIN(n7882),
    .SDIN_t(n7882_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7883),
    .Q_t(n7883_t),
    .QN(n6360),
    .QN_t(n6360_t)
  );


  sdffs1
  \DFF_1551/Q_reg 
  (
    .DIN(WX10858),
    .DIN_t(WX10858_t),
    .SDIN(n7881),
    .SDIN_t(n7881_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7882),
    .Q_t(n7882_t),
    .QN(n6361),
    .QN_t(n6361_t)
  );


  sdffs1
  \DFF_1550/Q_reg 
  (
    .DIN(WX10856),
    .DIN_t(WX10856_t),
    .SDIN(n7880),
    .SDIN_t(n7880_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7881),
    .Q_t(n7881_t),
    .QN(n6362),
    .QN_t(n6362_t)
  );


  sdffs1
  \DFF_1549/Q_reg 
  (
    .DIN(WX10854),
    .DIN_t(WX10854_t),
    .SDIN(n7879),
    .SDIN_t(n7879_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7880),
    .Q_t(n7880_t),
    .QN(n6363),
    .QN_t(n6363_t)
  );


  sdffs1
  \DFF_1548/Q_reg 
  (
    .DIN(WX10852),
    .DIN_t(WX10852_t),
    .SDIN(n7878),
    .SDIN_t(n7878_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7879),
    .Q_t(n7879_t),
    .QN(n6364),
    .QN_t(n6364_t)
  );


  sdffs1
  \DFF_1547/Q_reg 
  (
    .DIN(WX10850),
    .DIN_t(WX10850_t),
    .SDIN(n7877),
    .SDIN_t(n7877_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7878),
    .Q_t(n7878_t),
    .QN(n6365),
    .QN_t(n6365_t)
  );


  sdffs1
  \DFF_1546/Q_reg 
  (
    .DIN(WX10848),
    .DIN_t(WX10848_t),
    .SDIN(n7876),
    .SDIN_t(n7876_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7877),
    .Q_t(n7877_t),
    .QN(n6366),
    .QN_t(n6366_t)
  );


  sdffs1
  \DFF_1545/Q_reg 
  (
    .DIN(WX10846),
    .DIN_t(WX10846_t),
    .SDIN(n7875),
    .SDIN_t(n7875_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7876),
    .Q_t(n7876_t),
    .QN(n6367),
    .QN_t(n6367_t)
  );


  sdffs1
  \DFF_1544/Q_reg 
  (
    .DIN(WX10844),
    .DIN_t(WX10844_t),
    .SDIN(n7874),
    .SDIN_t(n7874_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7875),
    .Q_t(n7875_t),
    .QN(n6368),
    .QN_t(n6368_t)
  );


  sdffs1
  \DFF_1543/Q_reg 
  (
    .DIN(WX10842),
    .DIN_t(WX10842_t),
    .SDIN(n7873),
    .SDIN_t(n7873_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7874),
    .Q_t(n7874_t),
    .QN(n6369),
    .QN_t(n6369_t)
  );


  sdffs1
  \DFF_1542/Q_reg 
  (
    .DIN(WX10840),
    .DIN_t(WX10840_t),
    .SDIN(n7872),
    .SDIN_t(n7872_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7873),
    .Q_t(n7873_t),
    .QN(n6370),
    .QN_t(n6370_t)
  );


  sdffs1
  \DFF_1541/Q_reg 
  (
    .DIN(WX10838),
    .DIN_t(WX10838_t),
    .SDIN(n7871),
    .SDIN_t(n7871_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7872),
    .Q_t(n7872_t),
    .QN(n6371),
    .QN_t(n6371_t)
  );


  sdffs1
  \DFF_1540/Q_reg 
  (
    .DIN(WX10836),
    .DIN_t(WX10836_t),
    .SDIN(n7870),
    .SDIN_t(n7870_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7871),
    .Q_t(n7871_t),
    .QN(n6372),
    .QN_t(n6372_t)
  );


  sdffs1
  \DFF_1539/Q_reg 
  (
    .DIN(WX10834),
    .DIN_t(WX10834_t),
    .SDIN(n7869),
    .SDIN_t(n7869_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7870),
    .Q_t(n7870_t),
    .QN(n6373),
    .QN_t(n6373_t)
  );


  sdffs1
  \DFF_1538/Q_reg 
  (
    .DIN(WX10832),
    .DIN_t(WX10832_t),
    .SDIN(n7868),
    .SDIN_t(n7868_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7869),
    .Q_t(n7869_t),
    .QN(n6374),
    .QN_t(n6374_t)
  );


  sdffs1
  \DFF_1537/Q_reg 
  (
    .DIN(WX10830),
    .DIN_t(WX10830_t),
    .SDIN(n7867),
    .SDIN_t(n7867_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7868),
    .Q_t(n7868_t),
    .QN(n6375),
    .QN_t(n6375_t)
  );


  sdffs1
  \DFF_1536/Q_reg 
  (
    .DIN(WX10828),
    .DIN_t(WX10828_t),
    .SDIN(CRC_OUT_2_31),
    .SDIN_t(CRC_OUT_2_31_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7867),
    .Q_t(n7867_t),
    .QN(n6343),
    .QN_t(n6343_t)
  );


  sdffs1
  \DFF_1535/Q_reg 
  (
    .DIN(WX10377),
    .DIN_t(WX10377_t),
    .SDIN(CRC_OUT_2_30),
    .SDIN_t(CRC_OUT_2_30_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_31),
    .Q_t(CRC_OUT_2_31_t),
    .QN(n6430),
    .QN_t(n6430_t)
  );


  sdffs1
  \DFF_1534/Q_reg 
  (
    .DIN(WX10375),
    .DIN_t(WX10375_t),
    .SDIN(CRC_OUT_2_29),
    .SDIN_t(CRC_OUT_2_29_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_30),
    .Q_t(CRC_OUT_2_30_t),
    .QN(n6383),
    .QN_t(n6383_t)
  );


  sdffs1
  \DFF_1533/Q_reg 
  (
    .DIN(WX10373),
    .DIN_t(WX10373_t),
    .SDIN(CRC_OUT_2_28),
    .SDIN_t(CRC_OUT_2_28_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_29),
    .Q_t(CRC_OUT_2_29_t),
    .QN(n6385),
    .QN_t(n6385_t)
  );


  sdffs1
  \DFF_1532/Q_reg 
  (
    .DIN(WX10371),
    .DIN_t(WX10371_t),
    .SDIN(CRC_OUT_2_27),
    .SDIN_t(CRC_OUT_2_27_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_28),
    .Q_t(CRC_OUT_2_28_t),
    .QN(n6387),
    .QN_t(n6387_t)
  );


  sdffs1
  \DFF_1531/Q_reg 
  (
    .DIN(WX10369),
    .DIN_t(WX10369_t),
    .SDIN(CRC_OUT_2_26),
    .SDIN_t(CRC_OUT_2_26_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_27),
    .Q_t(CRC_OUT_2_27_t),
    .QN(n6389),
    .QN_t(n6389_t)
  );


  sdffs1
  \DFF_1530/Q_reg 
  (
    .DIN(WX10367),
    .DIN_t(WX10367_t),
    .SDIN(CRC_OUT_2_25),
    .SDIN_t(CRC_OUT_2_25_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_26),
    .Q_t(CRC_OUT_2_26_t),
    .QN(n6391),
    .QN_t(n6391_t)
  );


  sdffs1
  \DFF_1529/Q_reg 
  (
    .DIN(WX10365),
    .DIN_t(WX10365_t),
    .SDIN(CRC_OUT_2_24),
    .SDIN_t(CRC_OUT_2_24_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_25),
    .Q_t(CRC_OUT_2_25_t),
    .QN(n6393),
    .QN_t(n6393_t)
  );


  sdffs1
  \DFF_1528/Q_reg 
  (
    .DIN(WX10363),
    .DIN_t(WX10363_t),
    .SDIN(CRC_OUT_2_23),
    .SDIN_t(CRC_OUT_2_23_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_24),
    .Q_t(CRC_OUT_2_24_t),
    .QN(n6395),
    .QN_t(n6395_t)
  );


  sdffs1
  \DFF_1527/Q_reg 
  (
    .DIN(WX10361),
    .DIN_t(WX10361_t),
    .SDIN(CRC_OUT_2_22),
    .SDIN_t(CRC_OUT_2_22_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_23),
    .Q_t(CRC_OUT_2_23_t),
    .QN(n6397),
    .QN_t(n6397_t)
  );


  sdffs1
  \DFF_1526/Q_reg 
  (
    .DIN(WX10359),
    .DIN_t(WX10359_t),
    .SDIN(CRC_OUT_2_21),
    .SDIN_t(CRC_OUT_2_21_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_22),
    .Q_t(CRC_OUT_2_22_t),
    .QN(n6399),
    .QN_t(n6399_t)
  );


  sdffs1
  \DFF_1525/Q_reg 
  (
    .DIN(WX10357),
    .DIN_t(WX10357_t),
    .SDIN(CRC_OUT_2_20),
    .SDIN_t(CRC_OUT_2_20_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_21),
    .Q_t(CRC_OUT_2_21_t),
    .QN(n6401),
    .QN_t(n6401_t)
  );


  sdffs1
  \DFF_1524/Q_reg 
  (
    .DIN(WX10355),
    .DIN_t(WX10355_t),
    .SDIN(CRC_OUT_2_19),
    .SDIN_t(CRC_OUT_2_19_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_20),
    .Q_t(CRC_OUT_2_20_t),
    .QN(n6403),
    .QN_t(n6403_t)
  );


  sdffs1
  \DFF_1523/Q_reg 
  (
    .DIN(WX10353),
    .DIN_t(WX10353_t),
    .SDIN(CRC_OUT_2_18),
    .SDIN_t(CRC_OUT_2_18_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_19),
    .Q_t(CRC_OUT_2_19_t),
    .QN(n6405),
    .QN_t(n6405_t)
  );


  sdffs1
  \DFF_1522/Q_reg 
  (
    .DIN(WX10351),
    .DIN_t(WX10351_t),
    .SDIN(CRC_OUT_2_17),
    .SDIN_t(CRC_OUT_2_17_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_18),
    .Q_t(CRC_OUT_2_18_t),
    .QN(n6407),
    .QN_t(n6407_t)
  );


  sdffs1
  \DFF_1521/Q_reg 
  (
    .DIN(WX10349),
    .DIN_t(WX10349_t),
    .SDIN(CRC_OUT_2_16),
    .SDIN_t(CRC_OUT_2_16_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_17),
    .Q_t(CRC_OUT_2_17_t),
    .QN(n6409),
    .QN_t(n6409_t)
  );


  sdffs1
  \DFF_1520/Q_reg 
  (
    .DIN(WX10347),
    .DIN_t(WX10347_t),
    .SDIN(CRC_OUT_2_15),
    .SDIN_t(CRC_OUT_2_15_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_16),
    .Q_t(CRC_OUT_2_16_t),
    .QN(n6411),
    .QN_t(n6411_t)
  );


  sdffs1
  \DFF_1519/Q_reg 
  (
    .DIN(WX10345),
    .DIN_t(WX10345_t),
    .SDIN(CRC_OUT_2_14),
    .SDIN_t(CRC_OUT_2_14_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_15),
    .Q_t(CRC_OUT_2_15_t),
    .QN(n6413),
    .QN_t(n6413_t)
  );


  sdffs1
  \DFF_1518/Q_reg 
  (
    .DIN(WX10343),
    .DIN_t(WX10343_t),
    .SDIN(CRC_OUT_2_13),
    .SDIN_t(CRC_OUT_2_13_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_14),
    .Q_t(CRC_OUT_2_14_t),
    .QN(n6415),
    .QN_t(n6415_t)
  );


  sdffs1
  \DFF_1517/Q_reg 
  (
    .DIN(WX10341),
    .DIN_t(WX10341_t),
    .SDIN(CRC_OUT_2_12),
    .SDIN_t(CRC_OUT_2_12_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_13),
    .Q_t(CRC_OUT_2_13_t),
    .QN(n6416),
    .QN_t(n6416_t)
  );


  sdffs1
  \DFF_1516/Q_reg 
  (
    .DIN(WX10339),
    .DIN_t(WX10339_t),
    .SDIN(CRC_OUT_2_11),
    .SDIN_t(CRC_OUT_2_11_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_12),
    .Q_t(CRC_OUT_2_12_t),
    .QN(n6417),
    .QN_t(n6417_t)
  );


  sdffs1
  \DFF_1515/Q_reg 
  (
    .DIN(WX10337),
    .DIN_t(WX10337_t),
    .SDIN(CRC_OUT_2_10),
    .SDIN_t(CRC_OUT_2_10_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_11),
    .Q_t(CRC_OUT_2_11_t),
    .QN(n6418),
    .QN_t(n6418_t)
  );


  sdffs1
  \DFF_1514/Q_reg 
  (
    .DIN(WX10335),
    .DIN_t(WX10335_t),
    .SDIN(CRC_OUT_2_9),
    .SDIN_t(CRC_OUT_2_9_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_10),
    .Q_t(CRC_OUT_2_10_t),
    .QN(n6419),
    .QN_t(n6419_t)
  );


  sdffs1
  \DFF_1513/Q_reg 
  (
    .DIN(WX10333),
    .DIN_t(WX10333_t),
    .SDIN(CRC_OUT_2_8),
    .SDIN_t(CRC_OUT_2_8_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_9),
    .Q_t(CRC_OUT_2_9_t),
    .QN(n6420),
    .QN_t(n6420_t)
  );


  sdffs1
  \DFF_1512/Q_reg 
  (
    .DIN(WX10331),
    .DIN_t(WX10331_t),
    .SDIN(CRC_OUT_2_7),
    .SDIN_t(CRC_OUT_2_7_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_8),
    .Q_t(CRC_OUT_2_8_t),
    .QN(n6421),
    .QN_t(n6421_t)
  );


  sdffs1
  \DFF_1511/Q_reg 
  (
    .DIN(WX10329),
    .DIN_t(WX10329_t),
    .SDIN(CRC_OUT_2_6),
    .SDIN_t(CRC_OUT_2_6_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_7),
    .Q_t(CRC_OUT_2_7_t),
    .QN(n6422),
    .QN_t(n6422_t)
  );


  sdffs1
  \DFF_1510/Q_reg 
  (
    .DIN(WX10327),
    .DIN_t(WX10327_t),
    .SDIN(CRC_OUT_2_5),
    .SDIN_t(CRC_OUT_2_5_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_6),
    .Q_t(CRC_OUT_2_6_t),
    .QN(n6423),
    .QN_t(n6423_t)
  );


  sdffs1
  \DFF_1509/Q_reg 
  (
    .DIN(WX10325),
    .DIN_t(WX10325_t),
    .SDIN(CRC_OUT_2_4),
    .SDIN_t(CRC_OUT_2_4_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_5),
    .Q_t(CRC_OUT_2_5_t),
    .QN(n6424),
    .QN_t(n6424_t)
  );


  sdffs1
  \DFF_1508/Q_reg 
  (
    .DIN(WX10323),
    .DIN_t(WX10323_t),
    .SDIN(CRC_OUT_2_3),
    .SDIN_t(CRC_OUT_2_3_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_4),
    .Q_t(CRC_OUT_2_4_t),
    .QN(n6425),
    .QN_t(n6425_t)
  );


  sdffs1
  \DFF_1507/Q_reg 
  (
    .DIN(WX10321),
    .DIN_t(WX10321_t),
    .SDIN(CRC_OUT_2_2),
    .SDIN_t(CRC_OUT_2_2_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_3),
    .Q_t(CRC_OUT_2_3_t),
    .QN(n6426),
    .QN_t(n6426_t)
  );


  sdffs1
  \DFF_1506/Q_reg 
  (
    .DIN(WX10319),
    .DIN_t(WX10319_t),
    .SDIN(CRC_OUT_2_1),
    .SDIN_t(CRC_OUT_2_1_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_2),
    .Q_t(CRC_OUT_2_2_t),
    .QN(n6427),
    .QN_t(n6427_t)
  );


  sdffs1
  \DFF_1505/Q_reg 
  (
    .DIN(WX10317),
    .DIN_t(WX10317_t),
    .SDIN(CRC_OUT_2_0),
    .SDIN_t(CRC_OUT_2_0_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_1),
    .Q_t(CRC_OUT_2_1_t),
    .QN(n6428),
    .QN_t(n6428_t)
  );


  sdffs1
  \DFF_1504/Q_reg 
  (
    .DIN(WX10315),
    .DIN_t(WX10315_t),
    .SDIN(n7866),
    .SDIN_t(n7866_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_2_0),
    .Q_t(CRC_OUT_2_0_t),
    .QN(n6429),
    .QN_t(n6429_t)
  );


  sdffs1
  \DFF_1503/Q_reg 
  (
    .DIN(WX9949),
    .DIN_t(WX9949_t),
    .SDIN(n7865),
    .SDIN_t(n7865_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7866),
    .Q_t(n7866_t),
    .QN(n3205),
    .QN_t(n3205_t)
  );


  sdffs1
  \DFF_1502/Q_reg 
  (
    .DIN(WX9947),
    .DIN_t(WX9947_t),
    .SDIN(n7864),
    .SDIN_t(n7864_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7865),
    .Q_t(n7865_t),
    .QN(n3206),
    .QN_t(n3206_t)
  );


  sdffs1
  \DFF_1501/Q_reg 
  (
    .DIN(WX9945),
    .DIN_t(WX9945_t),
    .SDIN(n7863),
    .SDIN_t(n7863_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7864),
    .Q_t(n7864_t),
    .QN(n3207),
    .QN_t(n3207_t)
  );


  sdffs1
  \DFF_1500/Q_reg 
  (
    .DIN(WX9943),
    .DIN_t(WX9943_t),
    .SDIN(n7862),
    .SDIN_t(n7862_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7863),
    .Q_t(n7863_t),
    .QN(n3208),
    .QN_t(n3208_t)
  );


  sdffs1
  \DFF_1499/Q_reg 
  (
    .DIN(WX9941),
    .DIN_t(WX9941_t),
    .SDIN(n7861),
    .SDIN_t(n7861_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7862),
    .Q_t(n7862_t),
    .QN(n3209),
    .QN_t(n3209_t)
  );


  sdffs1
  \DFF_1498/Q_reg 
  (
    .DIN(WX9939),
    .DIN_t(WX9939_t),
    .SDIN(n7860),
    .SDIN_t(n7860_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7861),
    .Q_t(n7861_t),
    .QN(n3210),
    .QN_t(n3210_t)
  );


  sdffs1
  \DFF_1497/Q_reg 
  (
    .DIN(WX9937),
    .DIN_t(WX9937_t),
    .SDIN(n7859),
    .SDIN_t(n7859_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7860),
    .Q_t(n7860_t),
    .QN(n3211),
    .QN_t(n3211_t)
  );


  sdffs1
  \DFF_1496/Q_reg 
  (
    .DIN(WX9935),
    .DIN_t(WX9935_t),
    .SDIN(n7858),
    .SDIN_t(n7858_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7859),
    .Q_t(n7859_t),
    .QN(n3212),
    .QN_t(n3212_t)
  );


  sdffs1
  \DFF_1495/Q_reg 
  (
    .DIN(WX9933),
    .DIN_t(WX9933_t),
    .SDIN(n7857),
    .SDIN_t(n7857_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7858),
    .Q_t(n7858_t),
    .QN(n3213),
    .QN_t(n3213_t)
  );


  sdffs1
  \DFF_1494/Q_reg 
  (
    .DIN(WX9931),
    .DIN_t(WX9931_t),
    .SDIN(n7856),
    .SDIN_t(n7856_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7857),
    .Q_t(n7857_t),
    .QN(n3214),
    .QN_t(n3214_t)
  );


  sdffs1
  \DFF_1493/Q_reg 
  (
    .DIN(WX9929),
    .DIN_t(WX9929_t),
    .SDIN(n7855),
    .SDIN_t(n7855_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7856),
    .Q_t(n7856_t),
    .QN(n3215),
    .QN_t(n3215_t)
  );


  sdffs1
  \DFF_1492/Q_reg 
  (
    .DIN(WX9927),
    .DIN_t(WX9927_t),
    .SDIN(n7854),
    .SDIN_t(n7854_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7855),
    .Q_t(n7855_t),
    .QN(n3216),
    .QN_t(n3216_t)
  );


  sdffs1
  \DFF_1491/Q_reg 
  (
    .DIN(WX9925),
    .DIN_t(WX9925_t),
    .SDIN(n7853),
    .SDIN_t(n7853_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7854),
    .Q_t(n7854_t),
    .QN(n3217),
    .QN_t(n3217_t)
  );


  sdffs1
  \DFF_1490/Q_reg 
  (
    .DIN(WX9923),
    .DIN_t(WX9923_t),
    .SDIN(n7852),
    .SDIN_t(n7852_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7853),
    .Q_t(n7853_t),
    .QN(n3218),
    .QN_t(n3218_t)
  );


  sdffs1
  \DFF_1489/Q_reg 
  (
    .DIN(WX9921),
    .DIN_t(WX9921_t),
    .SDIN(n7851),
    .SDIN_t(n7851_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7852),
    .Q_t(n7852_t),
    .QN(n3219),
    .QN_t(n3219_t)
  );


  sdffs1
  \DFF_1488/Q_reg 
  (
    .DIN(WX9919),
    .DIN_t(WX9919_t),
    .SDIN(n7850),
    .SDIN_t(n7850_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7851),
    .Q_t(n7851_t),
    .QN(n3220),
    .QN_t(n3220_t)
  );


  sdffs1
  \DFF_1487/Q_reg 
  (
    .DIN(WX9917),
    .DIN_t(WX9917_t),
    .SDIN(n7849),
    .SDIN_t(n7849_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7850),
    .Q_t(n7850_t),
    .QN(n6414),
    .QN_t(n6414_t)
  );


  sdffs1
  \DFF_1486/Q_reg 
  (
    .DIN(WX9915),
    .DIN_t(WX9915_t),
    .SDIN(n7848),
    .SDIN_t(n7848_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7849),
    .Q_t(n7849_t),
    .QN(n6412),
    .QN_t(n6412_t)
  );


  sdffs1
  \DFF_1485/Q_reg 
  (
    .DIN(WX9913),
    .DIN_t(WX9913_t),
    .SDIN(n7847),
    .SDIN_t(n7847_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7848),
    .Q_t(n7848_t),
    .QN(n6410),
    .QN_t(n6410_t)
  );


  sdffs1
  \DFF_1484/Q_reg 
  (
    .DIN(WX9911),
    .DIN_t(WX9911_t),
    .SDIN(n7846),
    .SDIN_t(n7846_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7847),
    .Q_t(n7847_t),
    .QN(n6408),
    .QN_t(n6408_t)
  );


  sdffs1
  \DFF_1483/Q_reg 
  (
    .DIN(WX9909),
    .DIN_t(WX9909_t),
    .SDIN(n7845),
    .SDIN_t(n7845_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7846),
    .Q_t(n7846_t),
    .QN(n6406),
    .QN_t(n6406_t)
  );


  sdffs1
  \DFF_1482/Q_reg 
  (
    .DIN(WX9907),
    .DIN_t(WX9907_t),
    .SDIN(n7844),
    .SDIN_t(n7844_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7845),
    .Q_t(n7845_t),
    .QN(n6404),
    .QN_t(n6404_t)
  );


  sdffs1
  \DFF_1481/Q_reg 
  (
    .DIN(WX9905),
    .DIN_t(WX9905_t),
    .SDIN(n7843),
    .SDIN_t(n7843_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7844),
    .Q_t(n7844_t),
    .QN(n6402),
    .QN_t(n6402_t)
  );


  sdffs1
  \DFF_1480/Q_reg 
  (
    .DIN(WX9903),
    .DIN_t(WX9903_t),
    .SDIN(n7842),
    .SDIN_t(n7842_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7843),
    .Q_t(n7843_t),
    .QN(n6400),
    .QN_t(n6400_t)
  );


  sdffs1
  \DFF_1479/Q_reg 
  (
    .DIN(WX9901),
    .DIN_t(WX9901_t),
    .SDIN(n7841),
    .SDIN_t(n7841_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7842),
    .Q_t(n7842_t),
    .QN(n6398),
    .QN_t(n6398_t)
  );


  sdffs1
  \DFF_1478/Q_reg 
  (
    .DIN(WX9899),
    .DIN_t(WX9899_t),
    .SDIN(n7840),
    .SDIN_t(n7840_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7841),
    .Q_t(n7841_t),
    .QN(n6396),
    .QN_t(n6396_t)
  );


  sdffs1
  \DFF_1477/Q_reg 
  (
    .DIN(WX9897),
    .DIN_t(WX9897_t),
    .SDIN(n7839),
    .SDIN_t(n7839_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7840),
    .Q_t(n7840_t),
    .QN(n6394),
    .QN_t(n6394_t)
  );


  sdffs1
  \DFF_1476/Q_reg 
  (
    .DIN(WX9895),
    .DIN_t(WX9895_t),
    .SDIN(n7838),
    .SDIN_t(n7838_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7839),
    .Q_t(n7839_t),
    .QN(n6392),
    .QN_t(n6392_t)
  );


  sdffs1
  \DFF_1475/Q_reg 
  (
    .DIN(WX9893),
    .DIN_t(WX9893_t),
    .SDIN(n7837),
    .SDIN_t(n7837_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7838),
    .Q_t(n7838_t),
    .QN(n6390),
    .QN_t(n6390_t)
  );


  sdffs1
  \DFF_1474/Q_reg 
  (
    .DIN(WX9891),
    .DIN_t(WX9891_t),
    .SDIN(n7836),
    .SDIN_t(n7836_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7837),
    .Q_t(n7837_t),
    .QN(n6388),
    .QN_t(n6388_t)
  );


  sdffs1
  \DFF_1473/Q_reg 
  (
    .DIN(WX9889),
    .DIN_t(WX9889_t),
    .SDIN(n7835),
    .SDIN_t(n7835_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7836),
    .Q_t(n7836_t),
    .QN(n6386),
    .QN_t(n6386_t)
  );


  sdffs1
  \DFF_1472/Q_reg 
  (
    .DIN(WX9887),
    .DIN_t(WX9887_t),
    .SDIN(n7834),
    .SDIN_t(n7834_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7835),
    .Q_t(n7835_t),
    .QN(n6384),
    .QN_t(n6384_t)
  );


  sdffs1
  \DFF_1471/Q_reg 
  (
    .DIN(WX9885),
    .DIN_t(WX9885_t),
    .SDIN(n7833),
    .SDIN_t(n7833_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7834),
    .Q_t(n7834_t),
    .QN(n4997),
    .QN_t(n4997_t)
  );


  sdffs1
  \DFF_1470/Q_reg 
  (
    .DIN(WX9883),
    .DIN_t(WX9883_t),
    .SDIN(n7832),
    .SDIN_t(n7832_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7833),
    .Q_t(n7833_t),
    .QN(n5001),
    .QN_t(n5001_t)
  );


  sdffs1
  \DFF_1469/Q_reg 
  (
    .DIN(WX9881),
    .DIN_t(WX9881_t),
    .SDIN(n7831),
    .SDIN_t(n7831_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7832),
    .Q_t(n7832_t),
    .QN(n5005),
    .QN_t(n5005_t)
  );


  sdffs1
  \DFF_1468/Q_reg 
  (
    .DIN(WX9879),
    .DIN_t(WX9879_t),
    .SDIN(n7830),
    .SDIN_t(n7830_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7831),
    .Q_t(n7831_t),
    .QN(n5009),
    .QN_t(n5009_t)
  );


  sdffs1
  \DFF_1467/Q_reg 
  (
    .DIN(WX9877),
    .DIN_t(WX9877_t),
    .SDIN(n7829),
    .SDIN_t(n7829_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7830),
    .Q_t(n7830_t),
    .QN(n5013),
    .QN_t(n5013_t)
  );


  sdffs1
  \DFF_1466/Q_reg 
  (
    .DIN(WX9875),
    .DIN_t(WX9875_t),
    .SDIN(n7828),
    .SDIN_t(n7828_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7829),
    .Q_t(n7829_t),
    .QN(n5017),
    .QN_t(n5017_t)
  );


  sdffs1
  \DFF_1465/Q_reg 
  (
    .DIN(WX9873),
    .DIN_t(WX9873_t),
    .SDIN(n7827),
    .SDIN_t(n7827_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7828),
    .Q_t(n7828_t),
    .QN(n5021),
    .QN_t(n5021_t)
  );


  sdffs1
  \DFF_1464/Q_reg 
  (
    .DIN(WX9871),
    .DIN_t(WX9871_t),
    .SDIN(n7826),
    .SDIN_t(n7826_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7827),
    .Q_t(n7827_t),
    .QN(n5025),
    .QN_t(n5025_t)
  );


  sdffs1
  \DFF_1463/Q_reg 
  (
    .DIN(WX9869),
    .DIN_t(WX9869_t),
    .SDIN(n7825),
    .SDIN_t(n7825_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7826),
    .Q_t(n7826_t),
    .QN(n5029),
    .QN_t(n5029_t)
  );


  sdffs1
  \DFF_1462/Q_reg 
  (
    .DIN(WX9867),
    .DIN_t(WX9867_t),
    .SDIN(n7824),
    .SDIN_t(n7824_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7825),
    .Q_t(n7825_t),
    .QN(n5033),
    .QN_t(n5033_t)
  );


  sdffs1
  \DFF_1461/Q_reg 
  (
    .DIN(WX9865),
    .DIN_t(WX9865_t),
    .SDIN(n7823),
    .SDIN_t(n7823_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7824),
    .Q_t(n7824_t),
    .QN(n5037),
    .QN_t(n5037_t)
  );


  sdffs1
  \DFF_1460/Q_reg 
  (
    .DIN(WX9863),
    .DIN_t(WX9863_t),
    .SDIN(n7822),
    .SDIN_t(n7822_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7823),
    .Q_t(n7823_t),
    .QN(n5041),
    .QN_t(n5041_t)
  );


  sdffs1
  \DFF_1459/Q_reg 
  (
    .DIN(WX9861),
    .DIN_t(WX9861_t),
    .SDIN(n7821),
    .SDIN_t(n7821_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7822),
    .Q_t(n7822_t),
    .QN(n5045),
    .QN_t(n5045_t)
  );


  sdffs1
  \DFF_1458/Q_reg 
  (
    .DIN(WX9859),
    .DIN_t(WX9859_t),
    .SDIN(n7820),
    .SDIN_t(n7820_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7821),
    .Q_t(n7821_t),
    .QN(n5049),
    .QN_t(n5049_t)
  );


  sdffs1
  \DFF_1457/Q_reg 
  (
    .DIN(WX9857),
    .DIN_t(WX9857_t),
    .SDIN(n7819),
    .SDIN_t(n7819_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7820),
    .Q_t(n7820_t),
    .QN(n5053),
    .QN_t(n5053_t)
  );


  sdffs1
  \DFF_1456/Q_reg 
  (
    .DIN(WX9855),
    .DIN_t(WX9855_t),
    .SDIN(n7818),
    .SDIN_t(n7818_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7819),
    .Q_t(n7819_t),
    .QN(n5057),
    .QN_t(n5057_t)
  );


  sdffs1
  \DFF_1455/Q_reg 
  (
    .DIN(WX9853),
    .DIN_t(WX9853_t),
    .SDIN(n7817),
    .SDIN_t(n7817_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7818),
    .Q_t(n7818_t),
    .QN(n5061),
    .QN_t(n5061_t)
  );


  sdffs1
  \DFF_1454/Q_reg 
  (
    .DIN(WX9851),
    .DIN_t(WX9851_t),
    .SDIN(n7816),
    .SDIN_t(n7816_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7817),
    .Q_t(n7817_t),
    .QN(n5065),
    .QN_t(n5065_t)
  );


  sdffs1
  \DFF_1453/Q_reg 
  (
    .DIN(WX9849),
    .DIN_t(WX9849_t),
    .SDIN(n7815),
    .SDIN_t(n7815_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7816),
    .Q_t(n7816_t),
    .QN(n5069),
    .QN_t(n5069_t)
  );


  sdffs1
  \DFF_1452/Q_reg 
  (
    .DIN(WX9847),
    .DIN_t(WX9847_t),
    .SDIN(n7814),
    .SDIN_t(n7814_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7815),
    .Q_t(n7815_t),
    .QN(n5073),
    .QN_t(n5073_t)
  );


  sdffs1
  \DFF_1451/Q_reg 
  (
    .DIN(WX9845),
    .DIN_t(WX9845_t),
    .SDIN(n7813),
    .SDIN_t(n7813_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7814),
    .Q_t(n7814_t),
    .QN(n5077),
    .QN_t(n5077_t)
  );


  sdffs1
  \DFF_1450/Q_reg 
  (
    .DIN(WX9843),
    .DIN_t(WX9843_t),
    .SDIN(n7812),
    .SDIN_t(n7812_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7813),
    .Q_t(n7813_t),
    .QN(n5081),
    .QN_t(n5081_t)
  );


  sdffs1
  \DFF_1449/Q_reg 
  (
    .DIN(WX9841),
    .DIN_t(WX9841_t),
    .SDIN(n7811),
    .SDIN_t(n7811_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7812),
    .Q_t(n7812_t),
    .QN(n5085),
    .QN_t(n5085_t)
  );


  sdffs1
  \DFF_1448/Q_reg 
  (
    .DIN(WX9839),
    .DIN_t(WX9839_t),
    .SDIN(n7810),
    .SDIN_t(n7810_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7811),
    .Q_t(n7811_t),
    .QN(n5089),
    .QN_t(n5089_t)
  );


  sdffs1
  \DFF_1447/Q_reg 
  (
    .DIN(WX9837),
    .DIN_t(WX9837_t),
    .SDIN(n7809),
    .SDIN_t(n7809_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7810),
    .Q_t(n7810_t),
    .QN(n5093),
    .QN_t(n5093_t)
  );


  sdffs1
  \DFF_1446/Q_reg 
  (
    .DIN(WX9835),
    .DIN_t(WX9835_t),
    .SDIN(n7808),
    .SDIN_t(n7808_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7809),
    .Q_t(n7809_t),
    .QN(n5097),
    .QN_t(n5097_t)
  );


  sdffs1
  \DFF_1445/Q_reg 
  (
    .DIN(WX9833),
    .DIN_t(WX9833_t),
    .SDIN(n7807),
    .SDIN_t(n7807_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7808),
    .Q_t(n7808_t),
    .QN(n5101),
    .QN_t(n5101_t)
  );


  sdffs1
  \DFF_1444/Q_reg 
  (
    .DIN(WX9831),
    .DIN_t(WX9831_t),
    .SDIN(n7806),
    .SDIN_t(n7806_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7807),
    .Q_t(n7807_t),
    .QN(n5105),
    .QN_t(n5105_t)
  );


  sdffs1
  \DFF_1443/Q_reg 
  (
    .DIN(WX9829),
    .DIN_t(WX9829_t),
    .SDIN(n7805),
    .SDIN_t(n7805_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7806),
    .Q_t(n7806_t),
    .QN(n5109),
    .QN_t(n5109_t)
  );


  sdffs1
  \DFF_1442/Q_reg 
  (
    .DIN(WX9827),
    .DIN_t(WX9827_t),
    .SDIN(n7804),
    .SDIN_t(n7804_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7805),
    .Q_t(n7805_t),
    .QN(n5113),
    .QN_t(n5113_t)
  );


  sdffs1
  \DFF_1441/Q_reg 
  (
    .DIN(WX9825),
    .DIN_t(WX9825_t),
    .SDIN(n7803),
    .SDIN_t(n7803_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7804),
    .Q_t(n7804_t),
    .QN(n5117),
    .QN_t(n5117_t)
  );


  sdffs1
  \DFF_1440/Q_reg 
  (
    .DIN(WX9823),
    .DIN_t(WX9823_t),
    .SDIN(n7802),
    .SDIN_t(n7802_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7803),
    .Q_t(n7803_t),
    .QN(n5121),
    .QN_t(n5121_t)
  );


  sdffs1
  \DFF_1439/Q_reg 
  (
    .DIN(WX9821),
    .DIN_t(WX9821_t),
    .SDIN(n7801),
    .SDIN_t(n7801_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7802),
    .Q_t(n7802_t),
    .QN(n4996),
    .QN_t(n4996_t)
  );


  sdffs1
  \DFF_1438/Q_reg 
  (
    .DIN(WX9819),
    .DIN_t(WX9819_t),
    .SDIN(n7800),
    .SDIN_t(n7800_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7801),
    .Q_t(n7801_t),
    .QN(n5000),
    .QN_t(n5000_t)
  );


  sdffs1
  \DFF_1437/Q_reg 
  (
    .DIN(WX9817),
    .DIN_t(WX9817_t),
    .SDIN(n7799),
    .SDIN_t(n7799_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7800),
    .Q_t(n7800_t),
    .QN(n5004),
    .QN_t(n5004_t)
  );


  sdffs1
  \DFF_1436/Q_reg 
  (
    .DIN(WX9815),
    .DIN_t(WX9815_t),
    .SDIN(n7798),
    .SDIN_t(n7798_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7799),
    .Q_t(n7799_t),
    .QN(n5008),
    .QN_t(n5008_t)
  );


  sdffs1
  \DFF_1435/Q_reg 
  (
    .DIN(WX9813),
    .DIN_t(WX9813_t),
    .SDIN(n7797),
    .SDIN_t(n7797_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7798),
    .Q_t(n7798_t),
    .QN(n5012),
    .QN_t(n5012_t)
  );


  sdffs1
  \DFF_1434/Q_reg 
  (
    .DIN(WX9811),
    .DIN_t(WX9811_t),
    .SDIN(n7796),
    .SDIN_t(n7796_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7797),
    .Q_t(n7797_t),
    .QN(n5016),
    .QN_t(n5016_t)
  );


  sdffs1
  \DFF_1433/Q_reg 
  (
    .DIN(WX9809),
    .DIN_t(WX9809_t),
    .SDIN(n7795),
    .SDIN_t(n7795_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7796),
    .Q_t(n7796_t),
    .QN(n5020),
    .QN_t(n5020_t)
  );


  sdffs1
  \DFF_1432/Q_reg 
  (
    .DIN(WX9807),
    .DIN_t(WX9807_t),
    .SDIN(n7794),
    .SDIN_t(n7794_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7795),
    .Q_t(n7795_t),
    .QN(n5024),
    .QN_t(n5024_t)
  );


  sdffs1
  \DFF_1431/Q_reg 
  (
    .DIN(WX9805),
    .DIN_t(WX9805_t),
    .SDIN(n7793),
    .SDIN_t(n7793_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7794),
    .Q_t(n7794_t),
    .QN(n5028),
    .QN_t(n5028_t)
  );


  sdffs1
  \DFF_1430/Q_reg 
  (
    .DIN(WX9803),
    .DIN_t(WX9803_t),
    .SDIN(n7792),
    .SDIN_t(n7792_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7793),
    .Q_t(n7793_t),
    .QN(n5032),
    .QN_t(n5032_t)
  );


  sdffs1
  \DFF_1429/Q_reg 
  (
    .DIN(WX9801),
    .DIN_t(WX9801_t),
    .SDIN(n7791),
    .SDIN_t(n7791_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7792),
    .Q_t(n7792_t),
    .QN(n5036),
    .QN_t(n5036_t)
  );


  sdffs1
  \DFF_1428/Q_reg 
  (
    .DIN(WX9799),
    .DIN_t(WX9799_t),
    .SDIN(n7790),
    .SDIN_t(n7790_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7791),
    .Q_t(n7791_t),
    .QN(n5040),
    .QN_t(n5040_t)
  );


  sdffs1
  \DFF_1427/Q_reg 
  (
    .DIN(WX9797),
    .DIN_t(WX9797_t),
    .SDIN(n7789),
    .SDIN_t(n7789_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7790),
    .Q_t(n7790_t),
    .QN(n5044),
    .QN_t(n5044_t)
  );


  sdffs1
  \DFF_1426/Q_reg 
  (
    .DIN(WX9795),
    .DIN_t(WX9795_t),
    .SDIN(n7788),
    .SDIN_t(n7788_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7789),
    .Q_t(n7789_t),
    .QN(n5048),
    .QN_t(n5048_t)
  );


  sdffs1
  \DFF_1425/Q_reg 
  (
    .DIN(WX9793),
    .DIN_t(WX9793_t),
    .SDIN(n7787),
    .SDIN_t(n7787_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7788),
    .Q_t(n7788_t),
    .QN(n5052),
    .QN_t(n5052_t)
  );


  sdffs1
  \DFF_1424/Q_reg 
  (
    .DIN(WX9791),
    .DIN_t(WX9791_t),
    .SDIN(n5060),
    .SDIN_t(n5060_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7787),
    .Q_t(n7787_t),
    .QN(n5056),
    .QN_t(n5056_t)
  );


  sdffs1
  \DFF_1423/Q_reg 
  (
    .DIN(WX9789),
    .DIN_t(WX9789_t),
    .SDIN(n5064),
    .SDIN_t(n5064_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5060),
    .Q_t(n5060_t)
  );


  sdffs1
  \DFF_1422/Q_reg 
  (
    .DIN(WX9787),
    .DIN_t(WX9787_t),
    .SDIN(n5068),
    .SDIN_t(n5068_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5064),
    .Q_t(n5064_t)
  );


  sdffs1
  \DFF_1421/Q_reg 
  (
    .DIN(WX9785),
    .DIN_t(WX9785_t),
    .SDIN(n5072),
    .SDIN_t(n5072_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5068),
    .Q_t(n5068_t)
  );


  sdffs1
  \DFF_1420/Q_reg 
  (
    .DIN(WX9783),
    .DIN_t(WX9783_t),
    .SDIN(n5076),
    .SDIN_t(n5076_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5072),
    .Q_t(n5072_t)
  );


  sdffs1
  \DFF_1419/Q_reg 
  (
    .DIN(WX9781),
    .DIN_t(WX9781_t),
    .SDIN(n5080),
    .SDIN_t(n5080_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5076),
    .Q_t(n5076_t)
  );


  sdffs1
  \DFF_1418/Q_reg 
  (
    .DIN(WX9779),
    .DIN_t(WX9779_t),
    .SDIN(n5084),
    .SDIN_t(n5084_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5080),
    .Q_t(n5080_t)
  );


  sdffs1
  \DFF_1417/Q_reg 
  (
    .DIN(WX9777),
    .DIN_t(WX9777_t),
    .SDIN(n5088),
    .SDIN_t(n5088_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5084),
    .Q_t(n5084_t)
  );


  sdffs1
  \DFF_1416/Q_reg 
  (
    .DIN(WX9775),
    .DIN_t(WX9775_t),
    .SDIN(n5092),
    .SDIN_t(n5092_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5088),
    .Q_t(n5088_t)
  );


  sdffs1
  \DFF_1415/Q_reg 
  (
    .DIN(WX9773),
    .DIN_t(WX9773_t),
    .SDIN(n5096),
    .SDIN_t(n5096_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5092),
    .Q_t(n5092_t)
  );


  sdffs1
  \DFF_1414/Q_reg 
  (
    .DIN(WX9771),
    .DIN_t(WX9771_t),
    .SDIN(n5100),
    .SDIN_t(n5100_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5096),
    .Q_t(n5096_t)
  );


  sdffs1
  \DFF_1413/Q_reg 
  (
    .DIN(WX9769),
    .DIN_t(WX9769_t),
    .SDIN(n5104),
    .SDIN_t(n5104_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5100),
    .Q_t(n5100_t)
  );


  sdffs1
  \DFF_1412/Q_reg 
  (
    .DIN(WX9767),
    .DIN_t(WX9767_t),
    .SDIN(n5108),
    .SDIN_t(n5108_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5104),
    .Q_t(n5104_t)
  );


  sdffs1
  \DFF_1411/Q_reg 
  (
    .DIN(WX9765),
    .DIN_t(WX9765_t),
    .SDIN(n5112),
    .SDIN_t(n5112_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5108),
    .Q_t(n5108_t)
  );


  sdffs1
  \DFF_1410/Q_reg 
  (
    .DIN(WX9763),
    .DIN_t(WX9763_t),
    .SDIN(n5116),
    .SDIN_t(n5116_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5112),
    .Q_t(n5112_t)
  );


  sdffs1
  \DFF_1409/Q_reg 
  (
    .DIN(WX9761),
    .DIN_t(WX9761_t),
    .SDIN(n5120),
    .SDIN_t(n5120_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5116),
    .Q_t(n5116_t)
  );


  sdffs1
  \DFF_1408/Q_reg 
  (
    .DIN(WX9759),
    .DIN_t(WX9759_t),
    .SDIN(n4995),
    .SDIN_t(n4995_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5120),
    .Q_t(n5120_t)
  );


  sdffs1
  \DFF_1407/Q_reg 
  (
    .DIN(WX9757),
    .DIN_t(WX9757_t),
    .SDIN(n4999),
    .SDIN_t(n4999_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n4995),
    .Q_t(n4995_t)
  );


  sdffs1
  \DFF_1406/Q_reg 
  (
    .DIN(WX9755),
    .DIN_t(WX9755_t),
    .SDIN(n5003),
    .SDIN_t(n5003_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n4999),
    .Q_t(n4999_t)
  );


  sdffs1
  \DFF_1405/Q_reg 
  (
    .DIN(WX9753),
    .DIN_t(WX9753_t),
    .SDIN(n5007),
    .SDIN_t(n5007_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5003),
    .Q_t(n5003_t)
  );


  sdffs1
  \DFF_1404/Q_reg 
  (
    .DIN(WX9751),
    .DIN_t(WX9751_t),
    .SDIN(n5011),
    .SDIN_t(n5011_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5007),
    .Q_t(n5007_t)
  );


  sdffs1
  \DFF_1403/Q_reg 
  (
    .DIN(WX9749),
    .DIN_t(WX9749_t),
    .SDIN(n5015),
    .SDIN_t(n5015_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5011),
    .Q_t(n5011_t)
  );


  sdffs1
  \DFF_1402/Q_reg 
  (
    .DIN(WX9747),
    .DIN_t(WX9747_t),
    .SDIN(n5019),
    .SDIN_t(n5019_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5015),
    .Q_t(n5015_t)
  );


  sdffs1
  \DFF_1401/Q_reg 
  (
    .DIN(WX9745),
    .DIN_t(WX9745_t),
    .SDIN(n5023),
    .SDIN_t(n5023_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5019),
    .Q_t(n5019_t)
  );


  sdffs1
  \DFF_1400/Q_reg 
  (
    .DIN(WX9743),
    .DIN_t(WX9743_t),
    .SDIN(n5027),
    .SDIN_t(n5027_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5023),
    .Q_t(n5023_t)
  );


  sdffs1
  \DFF_1399/Q_reg 
  (
    .DIN(WX9741),
    .DIN_t(WX9741_t),
    .SDIN(n5031),
    .SDIN_t(n5031_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5027),
    .Q_t(n5027_t)
  );


  sdffs1
  \DFF_1398/Q_reg 
  (
    .DIN(WX9739),
    .DIN_t(WX9739_t),
    .SDIN(n5035),
    .SDIN_t(n5035_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5031),
    .Q_t(n5031_t)
  );


  sdffs1
  \DFF_1397/Q_reg 
  (
    .DIN(WX9737),
    .DIN_t(WX9737_t),
    .SDIN(n5039),
    .SDIN_t(n5039_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5035),
    .Q_t(n5035_t)
  );


  sdffs1
  \DFF_1396/Q_reg 
  (
    .DIN(WX9735),
    .DIN_t(WX9735_t),
    .SDIN(n5043),
    .SDIN_t(n5043_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5039),
    .Q_t(n5039_t)
  );


  sdffs1
  \DFF_1395/Q_reg 
  (
    .DIN(WX9733),
    .DIN_t(WX9733_t),
    .SDIN(n5047),
    .SDIN_t(n5047_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5043),
    .Q_t(n5043_t)
  );


  sdffs1
  \DFF_1394/Q_reg 
  (
    .DIN(WX9731),
    .DIN_t(WX9731_t),
    .SDIN(n5051),
    .SDIN_t(n5051_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5047),
    .Q_t(n5047_t)
  );


  sdffs1
  \DFF_1393/Q_reg 
  (
    .DIN(WX9729),
    .DIN_t(WX9729_t),
    .SDIN(n5055),
    .SDIN_t(n5055_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5051),
    .Q_t(n5051_t)
  );


  sdffs1
  \DFF_1392/Q_reg 
  (
    .DIN(WX9727),
    .DIN_t(WX9727_t),
    .SDIN(n7786),
    .SDIN_t(n7786_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5055),
    .Q_t(n5055_t)
  );


  sdffs1
  \DFF_1391/Q_reg 
  (
    .DIN(WX9725),
    .DIN_t(WX9725_t),
    .SDIN(n7785),
    .SDIN_t(n7785_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7786),
    .Q_t(n7786_t),
    .QN(n5059),
    .QN_t(n5059_t)
  );


  sdffs1
  \DFF_1390/Q_reg 
  (
    .DIN(WX9723),
    .DIN_t(WX9723_t),
    .SDIN(n7784),
    .SDIN_t(n7784_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7785),
    .Q_t(n7785_t),
    .QN(n5063),
    .QN_t(n5063_t)
  );


  sdffs1
  \DFF_1389/Q_reg 
  (
    .DIN(WX9721),
    .DIN_t(WX9721_t),
    .SDIN(n7783),
    .SDIN_t(n7783_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7784),
    .Q_t(n7784_t),
    .QN(n5067),
    .QN_t(n5067_t)
  );


  sdffs1
  \DFF_1388/Q_reg 
  (
    .DIN(WX9719),
    .DIN_t(WX9719_t),
    .SDIN(n7782),
    .SDIN_t(n7782_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7783),
    .Q_t(n7783_t),
    .QN(n5071),
    .QN_t(n5071_t)
  );


  sdffs1
  \DFF_1387/Q_reg 
  (
    .DIN(WX9717),
    .DIN_t(WX9717_t),
    .SDIN(n7781),
    .SDIN_t(n7781_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7782),
    .Q_t(n7782_t),
    .QN(n5075),
    .QN_t(n5075_t)
  );


  sdffs1
  \DFF_1386/Q_reg 
  (
    .DIN(WX9715),
    .DIN_t(WX9715_t),
    .SDIN(n7780),
    .SDIN_t(n7780_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7781),
    .Q_t(n7781_t),
    .QN(n5079),
    .QN_t(n5079_t)
  );


  sdffs1
  \DFF_1385/Q_reg 
  (
    .DIN(WX9713),
    .DIN_t(WX9713_t),
    .SDIN(n7779),
    .SDIN_t(n7779_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7780),
    .Q_t(n7780_t),
    .QN(n5083),
    .QN_t(n5083_t)
  );


  sdffs1
  \DFF_1384/Q_reg 
  (
    .DIN(WX9711),
    .DIN_t(WX9711_t),
    .SDIN(n7778),
    .SDIN_t(n7778_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7779),
    .Q_t(n7779_t),
    .QN(n5087),
    .QN_t(n5087_t)
  );


  sdffs1
  \DFF_1383/Q_reg 
  (
    .DIN(WX9709),
    .DIN_t(WX9709_t),
    .SDIN(n7777),
    .SDIN_t(n7777_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7778),
    .Q_t(n7778_t),
    .QN(n5091),
    .QN_t(n5091_t)
  );


  sdffs1
  \DFF_1382/Q_reg 
  (
    .DIN(WX9707),
    .DIN_t(WX9707_t),
    .SDIN(n7776),
    .SDIN_t(n7776_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7777),
    .Q_t(n7777_t),
    .QN(n5095),
    .QN_t(n5095_t)
  );


  sdffs1
  \DFF_1381/Q_reg 
  (
    .DIN(WX9705),
    .DIN_t(WX9705_t),
    .SDIN(n7775),
    .SDIN_t(n7775_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7776),
    .Q_t(n7776_t),
    .QN(n5099),
    .QN_t(n5099_t)
  );


  sdffs1
  \DFF_1380/Q_reg 
  (
    .DIN(WX9703),
    .DIN_t(WX9703_t),
    .SDIN(n7774),
    .SDIN_t(n7774_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7775),
    .Q_t(n7775_t),
    .QN(n5103),
    .QN_t(n5103_t)
  );


  sdffs1
  \DFF_1379/Q_reg 
  (
    .DIN(WX9701),
    .DIN_t(WX9701_t),
    .SDIN(n7773),
    .SDIN_t(n7773_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7774),
    .Q_t(n7774_t),
    .QN(n5107),
    .QN_t(n5107_t)
  );


  sdffs1
  \DFF_1378/Q_reg 
  (
    .DIN(WX9699),
    .DIN_t(WX9699_t),
    .SDIN(n7772),
    .SDIN_t(n7772_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7773),
    .Q_t(n7773_t),
    .QN(n5111),
    .QN_t(n5111_t)
  );


  sdffs1
  \DFF_1377/Q_reg 
  (
    .DIN(WX9697),
    .DIN_t(WX9697_t),
    .SDIN(n7771),
    .SDIN_t(n7771_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7772),
    .Q_t(n7772_t),
    .QN(n5115),
    .QN_t(n5115_t)
  );


  sdffs1
  \DFF_1376/Q_reg 
  (
    .DIN(WX9695),
    .DIN_t(WX9695_t),
    .SDIN(n7770),
    .SDIN_t(n7770_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7771),
    .Q_t(n7771_t),
    .QN(n5119),
    .QN_t(n5119_t)
  );


  sdffs1
  \DFF_1375/Q_reg 
  (
    .DIN(WX9597),
    .DIN_t(WX9597_t),
    .SDIN(n7769),
    .SDIN_t(n7769_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7770),
    .Q_t(n7770_t),
    .QN(n4964),
    .QN_t(n4964_t)
  );


  sdffs1
  \DFF_1374/Q_reg 
  (
    .DIN(WX9595),
    .DIN_t(WX9595_t),
    .SDIN(n7768),
    .SDIN_t(n7768_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7769),
    .Q_t(n7769_t),
    .QN(n4965),
    .QN_t(n4965_t)
  );


  sdffs1
  \DFF_1373/Q_reg 
  (
    .DIN(WX9593),
    .DIN_t(WX9593_t),
    .SDIN(n7767),
    .SDIN_t(n7767_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7768),
    .Q_t(n7768_t),
    .QN(n4966),
    .QN_t(n4966_t)
  );


  sdffs1
  \DFF_1372/Q_reg 
  (
    .DIN(WX9591),
    .DIN_t(WX9591_t),
    .SDIN(n7766),
    .SDIN_t(n7766_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7767),
    .Q_t(n7767_t),
    .QN(n4967),
    .QN_t(n4967_t)
  );


  sdffs1
  \DFF_1371/Q_reg 
  (
    .DIN(WX9589),
    .DIN_t(WX9589_t),
    .SDIN(n7765),
    .SDIN_t(n7765_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7766),
    .Q_t(n7766_t),
    .QN(n4968),
    .QN_t(n4968_t)
  );


  sdffs1
  \DFF_1370/Q_reg 
  (
    .DIN(WX9587),
    .DIN_t(WX9587_t),
    .SDIN(n7764),
    .SDIN_t(n7764_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7765),
    .Q_t(n7765_t),
    .QN(n4969),
    .QN_t(n4969_t)
  );


  sdffs1
  \DFF_1369/Q_reg 
  (
    .DIN(WX9585),
    .DIN_t(WX9585_t),
    .SDIN(n7763),
    .SDIN_t(n7763_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7764),
    .Q_t(n7764_t),
    .QN(n4970),
    .QN_t(n4970_t)
  );


  sdffs1
  \DFF_1368/Q_reg 
  (
    .DIN(WX9583),
    .DIN_t(WX9583_t),
    .SDIN(n7762),
    .SDIN_t(n7762_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7763),
    .Q_t(n7763_t),
    .QN(n4971),
    .QN_t(n4971_t)
  );


  sdffs1
  \DFF_1367/Q_reg 
  (
    .DIN(WX9581),
    .DIN_t(WX9581_t),
    .SDIN(n7761),
    .SDIN_t(n7761_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7762),
    .Q_t(n7762_t),
    .QN(n4972),
    .QN_t(n4972_t)
  );


  sdffs1
  \DFF_1366/Q_reg 
  (
    .DIN(WX9579),
    .DIN_t(WX9579_t),
    .SDIN(n7760),
    .SDIN_t(n7760_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7761),
    .Q_t(n7761_t),
    .QN(n4973),
    .QN_t(n4973_t)
  );


  sdffs1
  \DFF_1365/Q_reg 
  (
    .DIN(WX9577),
    .DIN_t(WX9577_t),
    .SDIN(n7759),
    .SDIN_t(n7759_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7760),
    .Q_t(n7760_t),
    .QN(n4974),
    .QN_t(n4974_t)
  );


  sdffs1
  \DFF_1364/Q_reg 
  (
    .DIN(WX9575),
    .DIN_t(WX9575_t),
    .SDIN(n7758),
    .SDIN_t(n7758_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7759),
    .Q_t(n7759_t),
    .QN(n4975),
    .QN_t(n4975_t)
  );


  sdffs1
  \DFF_1363/Q_reg 
  (
    .DIN(WX9573),
    .DIN_t(WX9573_t),
    .SDIN(n7757),
    .SDIN_t(n7757_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7758),
    .Q_t(n7758_t),
    .QN(n4976),
    .QN_t(n4976_t)
  );


  sdffs1
  \DFF_1362/Q_reg 
  (
    .DIN(WX9571),
    .DIN_t(WX9571_t),
    .SDIN(n7756),
    .SDIN_t(n7756_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7757),
    .Q_t(n7757_t),
    .QN(n4977),
    .QN_t(n4977_t)
  );


  sdffs1
  \DFF_1361/Q_reg 
  (
    .DIN(WX9569),
    .DIN_t(WX9569_t),
    .SDIN(n7755),
    .SDIN_t(n7755_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7756),
    .Q_t(n7756_t),
    .QN(n4978),
    .QN_t(n4978_t)
  );


  sdffs1
  \DFF_1360/Q_reg 
  (
    .DIN(WX9567),
    .DIN_t(WX9567_t),
    .SDIN(n7754),
    .SDIN_t(n7754_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7755),
    .Q_t(n7755_t),
    .QN(n4979),
    .QN_t(n4979_t)
  );


  sdffs1
  \DFF_1359/Q_reg 
  (
    .DIN(WX9565),
    .DIN_t(WX9565_t),
    .SDIN(n7753),
    .SDIN_t(n7753_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7754),
    .Q_t(n7754_t),
    .QN(n4980),
    .QN_t(n4980_t)
  );


  sdffs1
  \DFF_1358/Q_reg 
  (
    .DIN(WX9563),
    .DIN_t(WX9563_t),
    .SDIN(n7752),
    .SDIN_t(n7752_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7753),
    .Q_t(n7753_t),
    .QN(n4981),
    .QN_t(n4981_t)
  );


  sdffs1
  \DFF_1357/Q_reg 
  (
    .DIN(WX9561),
    .DIN_t(WX9561_t),
    .SDIN(n7751),
    .SDIN_t(n7751_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7752),
    .Q_t(n7752_t),
    .QN(n4982),
    .QN_t(n4982_t)
  );


  sdffs1
  \DFF_1356/Q_reg 
  (
    .DIN(WX9559),
    .DIN_t(WX9559_t),
    .SDIN(n7750),
    .SDIN_t(n7750_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7751),
    .Q_t(n7751_t),
    .QN(n4983),
    .QN_t(n4983_t)
  );


  sdffs1
  \DFF_1355/Q_reg 
  (
    .DIN(WX9557),
    .DIN_t(WX9557_t),
    .SDIN(n7749),
    .SDIN_t(n7749_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7750),
    .Q_t(n7750_t),
    .QN(n4984),
    .QN_t(n4984_t)
  );


  sdffs1
  \DFF_1354/Q_reg 
  (
    .DIN(WX9555),
    .DIN_t(WX9555_t),
    .SDIN(n7748),
    .SDIN_t(n7748_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7749),
    .Q_t(n7749_t),
    .QN(n4985),
    .QN_t(n4985_t)
  );


  sdffs1
  \DFF_1353/Q_reg 
  (
    .DIN(WX9553),
    .DIN_t(WX9553_t),
    .SDIN(n7747),
    .SDIN_t(n7747_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7748),
    .Q_t(n7748_t),
    .QN(n4986),
    .QN_t(n4986_t)
  );


  sdffs1
  \DFF_1352/Q_reg 
  (
    .DIN(WX9551),
    .DIN_t(WX9551_t),
    .SDIN(n7746),
    .SDIN_t(n7746_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7747),
    .Q_t(n7747_t),
    .QN(n4987),
    .QN_t(n4987_t)
  );


  sdffs1
  \DFF_1351/Q_reg 
  (
    .DIN(WX9549),
    .DIN_t(WX9549_t),
    .SDIN(n7745),
    .SDIN_t(n7745_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7746),
    .Q_t(n7746_t),
    .QN(n4988),
    .QN_t(n4988_t)
  );


  sdffs1
  \DFF_1350/Q_reg 
  (
    .DIN(WX9547),
    .DIN_t(WX9547_t),
    .SDIN(n7744),
    .SDIN_t(n7744_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7745),
    .Q_t(n7745_t),
    .QN(n4989),
    .QN_t(n4989_t)
  );


  sdffs1
  \DFF_1349/Q_reg 
  (
    .DIN(WX9545),
    .DIN_t(WX9545_t),
    .SDIN(n7743),
    .SDIN_t(n7743_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7744),
    .Q_t(n7744_t),
    .QN(n4990),
    .QN_t(n4990_t)
  );


  sdffs1
  \DFF_1348/Q_reg 
  (
    .DIN(WX9543),
    .DIN_t(WX9543_t),
    .SDIN(n7742),
    .SDIN_t(n7742_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7743),
    .Q_t(n7743_t),
    .QN(n4991),
    .QN_t(n4991_t)
  );


  sdffs1
  \DFF_1347/Q_reg 
  (
    .DIN(WX9541),
    .DIN_t(WX9541_t),
    .SDIN(n7741),
    .SDIN_t(n7741_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7742),
    .Q_t(n7742_t),
    .QN(n4992),
    .QN_t(n4992_t)
  );


  sdffs1
  \DFF_1346/Q_reg 
  (
    .DIN(WX9539),
    .DIN_t(WX9539_t),
    .SDIN(n7740),
    .SDIN_t(n7740_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7741),
    .Q_t(n7741_t),
    .QN(n4993),
    .QN_t(n4993_t)
  );


  sdffs1
  \DFF_1345/Q_reg 
  (
    .DIN(WX9537),
    .DIN_t(WX9537_t),
    .SDIN(n7739),
    .SDIN_t(n7739_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7740),
    .Q_t(n7740_t),
    .QN(n4994),
    .QN_t(n4994_t)
  );


  sdffs1
  \DFF_1344/Q_reg 
  (
    .DIN(WX9535),
    .DIN_t(WX9535_t),
    .SDIN(CRC_OUT_3_31),
    .SDIN_t(CRC_OUT_3_31_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7739),
    .Q_t(n7739_t),
    .QN(n4963),
    .QN_t(n4963_t)
  );


  sdffs1
  \DFF_1343/Q_reg 
  (
    .DIN(WX9084),
    .DIN_t(WX9084_t),
    .SDIN(CRC_OUT_3_30),
    .SDIN_t(CRC_OUT_3_30_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_31),
    .Q_t(CRC_OUT_3_31_t),
    .QN(n5122),
    .QN_t(n5122_t)
  );


  sdffs1
  \DFF_1342/Q_reg 
  (
    .DIN(WX9082),
    .DIN_t(WX9082_t),
    .SDIN(CRC_OUT_3_29),
    .SDIN_t(CRC_OUT_3_29_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_30),
    .Q_t(CRC_OUT_3_30_t),
    .QN(n5118),
    .QN_t(n5118_t)
  );


  sdffs1
  \DFF_1341/Q_reg 
  (
    .DIN(WX9080),
    .DIN_t(WX9080_t),
    .SDIN(CRC_OUT_3_28),
    .SDIN_t(CRC_OUT_3_28_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_29),
    .Q_t(CRC_OUT_3_29_t),
    .QN(n5114),
    .QN_t(n5114_t)
  );


  sdffs1
  \DFF_1340/Q_reg 
  (
    .DIN(WX9078),
    .DIN_t(WX9078_t),
    .SDIN(CRC_OUT_3_27),
    .SDIN_t(CRC_OUT_3_27_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_28),
    .Q_t(CRC_OUT_3_28_t),
    .QN(n5110),
    .QN_t(n5110_t)
  );


  sdffs1
  \DFF_1339/Q_reg 
  (
    .DIN(WX9076),
    .DIN_t(WX9076_t),
    .SDIN(CRC_OUT_3_26),
    .SDIN_t(CRC_OUT_3_26_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_27),
    .Q_t(CRC_OUT_3_27_t),
    .QN(n5106),
    .QN_t(n5106_t)
  );


  sdffs1
  \DFF_1338/Q_reg 
  (
    .DIN(WX9074),
    .DIN_t(WX9074_t),
    .SDIN(CRC_OUT_3_25),
    .SDIN_t(CRC_OUT_3_25_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_26),
    .Q_t(CRC_OUT_3_26_t),
    .QN(n5102),
    .QN_t(n5102_t)
  );


  sdffs1
  \DFF_1337/Q_reg 
  (
    .DIN(WX9072),
    .DIN_t(WX9072_t),
    .SDIN(CRC_OUT_3_24),
    .SDIN_t(CRC_OUT_3_24_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_25),
    .Q_t(CRC_OUT_3_25_t),
    .QN(n5098),
    .QN_t(n5098_t)
  );


  sdffs1
  \DFF_1336/Q_reg 
  (
    .DIN(WX9070),
    .DIN_t(WX9070_t),
    .SDIN(CRC_OUT_3_23),
    .SDIN_t(CRC_OUT_3_23_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_24),
    .Q_t(CRC_OUT_3_24_t),
    .QN(n5094),
    .QN_t(n5094_t)
  );


  sdffs1
  \DFF_1335/Q_reg 
  (
    .DIN(WX9068),
    .DIN_t(WX9068_t),
    .SDIN(CRC_OUT_3_22),
    .SDIN_t(CRC_OUT_3_22_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_23),
    .Q_t(CRC_OUT_3_23_t),
    .QN(n5090),
    .QN_t(n5090_t)
  );


  sdffs1
  \DFF_1334/Q_reg 
  (
    .DIN(WX9066),
    .DIN_t(WX9066_t),
    .SDIN(CRC_OUT_3_21),
    .SDIN_t(CRC_OUT_3_21_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_22),
    .Q_t(CRC_OUT_3_22_t),
    .QN(n5086),
    .QN_t(n5086_t)
  );


  sdffs1
  \DFF_1333/Q_reg 
  (
    .DIN(WX9064),
    .DIN_t(WX9064_t),
    .SDIN(CRC_OUT_3_20),
    .SDIN_t(CRC_OUT_3_20_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_21),
    .Q_t(CRC_OUT_3_21_t),
    .QN(n5082),
    .QN_t(n5082_t)
  );


  sdffs1
  \DFF_1332/Q_reg 
  (
    .DIN(WX9062),
    .DIN_t(WX9062_t),
    .SDIN(CRC_OUT_3_19),
    .SDIN_t(CRC_OUT_3_19_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_20),
    .Q_t(CRC_OUT_3_20_t),
    .QN(n5078),
    .QN_t(n5078_t)
  );


  sdffs1
  \DFF_1331/Q_reg 
  (
    .DIN(WX9060),
    .DIN_t(WX9060_t),
    .SDIN(CRC_OUT_3_18),
    .SDIN_t(CRC_OUT_3_18_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_19),
    .Q_t(CRC_OUT_3_19_t),
    .QN(n5074),
    .QN_t(n5074_t)
  );


  sdffs1
  \DFF_1330/Q_reg 
  (
    .DIN(WX9058),
    .DIN_t(WX9058_t),
    .SDIN(CRC_OUT_3_17),
    .SDIN_t(CRC_OUT_3_17_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_18),
    .Q_t(CRC_OUT_3_18_t),
    .QN(n5070),
    .QN_t(n5070_t)
  );


  sdffs1
  \DFF_1329/Q_reg 
  (
    .DIN(WX9056),
    .DIN_t(WX9056_t),
    .SDIN(CRC_OUT_3_16),
    .SDIN_t(CRC_OUT_3_16_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_17),
    .Q_t(CRC_OUT_3_17_t),
    .QN(n5066),
    .QN_t(n5066_t)
  );


  sdffs1
  \DFF_1328/Q_reg 
  (
    .DIN(WX9054),
    .DIN_t(WX9054_t),
    .SDIN(CRC_OUT_3_15),
    .SDIN_t(CRC_OUT_3_15_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_16),
    .Q_t(CRC_OUT_3_16_t),
    .QN(n5062),
    .QN_t(n5062_t)
  );


  sdffs1
  \DFF_1327/Q_reg 
  (
    .DIN(WX9052),
    .DIN_t(WX9052_t),
    .SDIN(CRC_OUT_3_14),
    .SDIN_t(CRC_OUT_3_14_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_15),
    .Q_t(CRC_OUT_3_15_t),
    .QN(n5058),
    .QN_t(n5058_t)
  );


  sdffs1
  \DFF_1326/Q_reg 
  (
    .DIN(WX9050),
    .DIN_t(WX9050_t),
    .SDIN(CRC_OUT_3_13),
    .SDIN_t(CRC_OUT_3_13_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_14),
    .Q_t(CRC_OUT_3_14_t),
    .QN(n5054),
    .QN_t(n5054_t)
  );


  sdffs1
  \DFF_1325/Q_reg 
  (
    .DIN(WX9048),
    .DIN_t(WX9048_t),
    .SDIN(CRC_OUT_3_12),
    .SDIN_t(CRC_OUT_3_12_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_13),
    .Q_t(CRC_OUT_3_13_t),
    .QN(n5050),
    .QN_t(n5050_t)
  );


  sdffs1
  \DFF_1324/Q_reg 
  (
    .DIN(WX9046),
    .DIN_t(WX9046_t),
    .SDIN(CRC_OUT_3_11),
    .SDIN_t(CRC_OUT_3_11_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_12),
    .Q_t(CRC_OUT_3_12_t),
    .QN(n5046),
    .QN_t(n5046_t)
  );


  sdffs1
  \DFF_1323/Q_reg 
  (
    .DIN(WX9044),
    .DIN_t(WX9044_t),
    .SDIN(CRC_OUT_3_10),
    .SDIN_t(CRC_OUT_3_10_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_11),
    .Q_t(CRC_OUT_3_11_t),
    .QN(n5042),
    .QN_t(n5042_t)
  );


  sdffs1
  \DFF_1322/Q_reg 
  (
    .DIN(WX9042),
    .DIN_t(WX9042_t),
    .SDIN(CRC_OUT_3_9),
    .SDIN_t(CRC_OUT_3_9_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_10),
    .Q_t(CRC_OUT_3_10_t),
    .QN(n5038),
    .QN_t(n5038_t)
  );


  sdffs1
  \DFF_1321/Q_reg 
  (
    .DIN(WX9040),
    .DIN_t(WX9040_t),
    .SDIN(CRC_OUT_3_8),
    .SDIN_t(CRC_OUT_3_8_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_9),
    .Q_t(CRC_OUT_3_9_t),
    .QN(n5034),
    .QN_t(n5034_t)
  );


  sdffs1
  \DFF_1320/Q_reg 
  (
    .DIN(WX9038),
    .DIN_t(WX9038_t),
    .SDIN(CRC_OUT_3_7),
    .SDIN_t(CRC_OUT_3_7_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_8),
    .Q_t(CRC_OUT_3_8_t),
    .QN(n5030),
    .QN_t(n5030_t)
  );


  sdffs1
  \DFF_1319/Q_reg 
  (
    .DIN(WX9036),
    .DIN_t(WX9036_t),
    .SDIN(CRC_OUT_3_6),
    .SDIN_t(CRC_OUT_3_6_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_7),
    .Q_t(CRC_OUT_3_7_t),
    .QN(n5026),
    .QN_t(n5026_t)
  );


  sdffs1
  \DFF_1318/Q_reg 
  (
    .DIN(WX9034),
    .DIN_t(WX9034_t),
    .SDIN(CRC_OUT_3_5),
    .SDIN_t(CRC_OUT_3_5_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_6),
    .Q_t(CRC_OUT_3_6_t),
    .QN(n5022),
    .QN_t(n5022_t)
  );


  sdffs1
  \DFF_1317/Q_reg 
  (
    .DIN(WX9032),
    .DIN_t(WX9032_t),
    .SDIN(CRC_OUT_3_4),
    .SDIN_t(CRC_OUT_3_4_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_5),
    .Q_t(CRC_OUT_3_5_t),
    .QN(n5018),
    .QN_t(n5018_t)
  );


  sdffs1
  \DFF_1316/Q_reg 
  (
    .DIN(WX9030),
    .DIN_t(WX9030_t),
    .SDIN(CRC_OUT_3_3),
    .SDIN_t(CRC_OUT_3_3_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_4),
    .Q_t(CRC_OUT_3_4_t),
    .QN(n5014),
    .QN_t(n5014_t)
  );


  sdffs1
  \DFF_1315/Q_reg 
  (
    .DIN(WX9028),
    .DIN_t(WX9028_t),
    .SDIN(CRC_OUT_3_2),
    .SDIN_t(CRC_OUT_3_2_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_3),
    .Q_t(CRC_OUT_3_3_t),
    .QN(n5010),
    .QN_t(n5010_t)
  );


  sdffs1
  \DFF_1314/Q_reg 
  (
    .DIN(WX9026),
    .DIN_t(WX9026_t),
    .SDIN(CRC_OUT_3_1),
    .SDIN_t(CRC_OUT_3_1_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_2),
    .Q_t(CRC_OUT_3_2_t),
    .QN(n5006),
    .QN_t(n5006_t)
  );


  sdffs1
  \DFF_1313/Q_reg 
  (
    .DIN(WX9024),
    .DIN_t(WX9024_t),
    .SDIN(CRC_OUT_3_0),
    .SDIN_t(CRC_OUT_3_0_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_1),
    .Q_t(CRC_OUT_3_1_t),
    .QN(n5002),
    .QN_t(n5002_t)
  );


  sdffs1
  \DFF_1312/Q_reg 
  (
    .DIN(WX9022),
    .DIN_t(WX9022_t),
    .SDIN(n7738),
    .SDIN_t(n7738_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_3_0),
    .Q_t(CRC_OUT_3_0_t),
    .QN(n4998),
    .QN_t(n4998_t)
  );


  sdffs1
  \DFF_1311/Q_reg 
  (
    .DIN(WX8656),
    .DIN_t(WX8656_t),
    .SDIN(n7737),
    .SDIN_t(n7737_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7738),
    .Q_t(n7738_t),
    .QN(n3221),
    .QN_t(n3221_t)
  );


  sdffs1
  \DFF_1310/Q_reg 
  (
    .DIN(WX8654),
    .DIN_t(WX8654_t),
    .SDIN(n7736),
    .SDIN_t(n7736_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7737),
    .Q_t(n7737_t),
    .QN(n3222),
    .QN_t(n3222_t)
  );


  sdffs1
  \DFF_1309/Q_reg 
  (
    .DIN(WX8652),
    .DIN_t(WX8652_t),
    .SDIN(n7735),
    .SDIN_t(n7735_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7736),
    .Q_t(n7736_t),
    .QN(n3223),
    .QN_t(n3223_t)
  );


  sdffs1
  \DFF_1308/Q_reg 
  (
    .DIN(WX8650),
    .DIN_t(WX8650_t),
    .SDIN(n7734),
    .SDIN_t(n7734_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7735),
    .Q_t(n7735_t),
    .QN(n3224),
    .QN_t(n3224_t)
  );


  sdffs1
  \DFF_1307/Q_reg 
  (
    .DIN(WX8648),
    .DIN_t(WX8648_t),
    .SDIN(n7733),
    .SDIN_t(n7733_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7734),
    .Q_t(n7734_t),
    .QN(n3225),
    .QN_t(n3225_t)
  );


  sdffs1
  \DFF_1306/Q_reg 
  (
    .DIN(WX8646),
    .DIN_t(WX8646_t),
    .SDIN(n7732),
    .SDIN_t(n7732_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7733),
    .Q_t(n7733_t),
    .QN(n3226),
    .QN_t(n3226_t)
  );


  sdffs1
  \DFF_1305/Q_reg 
  (
    .DIN(WX8644),
    .DIN_t(WX8644_t),
    .SDIN(n7731),
    .SDIN_t(n7731_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7732),
    .Q_t(n7732_t),
    .QN(n3227),
    .QN_t(n3227_t)
  );


  sdffs1
  \DFF_1304/Q_reg 
  (
    .DIN(WX8642),
    .DIN_t(WX8642_t),
    .SDIN(n7730),
    .SDIN_t(n7730_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7731),
    .Q_t(n7731_t),
    .QN(n3228),
    .QN_t(n3228_t)
  );


  sdffs1
  \DFF_1303/Q_reg 
  (
    .DIN(WX8640),
    .DIN_t(WX8640_t),
    .SDIN(n7729),
    .SDIN_t(n7729_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7730),
    .Q_t(n7730_t),
    .QN(n3229),
    .QN_t(n3229_t)
  );


  sdffs1
  \DFF_1302/Q_reg 
  (
    .DIN(WX8638),
    .DIN_t(WX8638_t),
    .SDIN(n7728),
    .SDIN_t(n7728_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7729),
    .Q_t(n7729_t),
    .QN(n3230),
    .QN_t(n3230_t)
  );


  sdffs1
  \DFF_1301/Q_reg 
  (
    .DIN(WX8636),
    .DIN_t(WX8636_t),
    .SDIN(n7727),
    .SDIN_t(n7727_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7728),
    .Q_t(n7728_t),
    .QN(n3231),
    .QN_t(n3231_t)
  );


  sdffs1
  \DFF_1300/Q_reg 
  (
    .DIN(WX8634),
    .DIN_t(WX8634_t),
    .SDIN(n7726),
    .SDIN_t(n7726_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7727),
    .Q_t(n7727_t),
    .QN(n3232),
    .QN_t(n3232_t)
  );


  sdffs1
  \DFF_1299/Q_reg 
  (
    .DIN(WX8632),
    .DIN_t(WX8632_t),
    .SDIN(n7725),
    .SDIN_t(n7725_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7726),
    .Q_t(n7726_t),
    .QN(n3233),
    .QN_t(n3233_t)
  );


  sdffs1
  \DFF_1298/Q_reg 
  (
    .DIN(WX8630),
    .DIN_t(WX8630_t),
    .SDIN(n7724),
    .SDIN_t(n7724_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7725),
    .Q_t(n7725_t),
    .QN(n3234),
    .QN_t(n3234_t)
  );


  sdffs1
  \DFF_1297/Q_reg 
  (
    .DIN(WX8628),
    .DIN_t(WX8628_t),
    .SDIN(n7723),
    .SDIN_t(n7723_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7724),
    .Q_t(n7724_t),
    .QN(n3235),
    .QN_t(n3235_t)
  );


  sdffs1
  \DFF_1296/Q_reg 
  (
    .DIN(WX8626),
    .DIN_t(WX8626_t),
    .SDIN(n7722),
    .SDIN_t(n7722_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7723),
    .Q_t(n7723_t),
    .QN(n3236),
    .QN_t(n3236_t)
  );


  sdffs1
  \DFF_1295/Q_reg 
  (
    .DIN(WX8624),
    .DIN_t(WX8624_t),
    .SDIN(n7721),
    .SDIN_t(n7721_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7722),
    .Q_t(n7722_t),
    .QN(n5222),
    .QN_t(n5222_t)
  );


  sdffs1
  \DFF_1294/Q_reg 
  (
    .DIN(WX8622),
    .DIN_t(WX8622_t),
    .SDIN(n7720),
    .SDIN_t(n7720_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7721),
    .Q_t(n7721_t),
    .QN(n5227),
    .QN_t(n5227_t)
  );


  sdffs1
  \DFF_1293/Q_reg 
  (
    .DIN(WX8620),
    .DIN_t(WX8620_t),
    .SDIN(n7719),
    .SDIN_t(n7719_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7720),
    .Q_t(n7720_t),
    .QN(n5232),
    .QN_t(n5232_t)
  );


  sdffs1
  \DFF_1292/Q_reg 
  (
    .DIN(WX8618),
    .DIN_t(WX8618_t),
    .SDIN(n7718),
    .SDIN_t(n7718_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7719),
    .Q_t(n7719_t),
    .QN(n5237),
    .QN_t(n5237_t)
  );


  sdffs1
  \DFF_1291/Q_reg 
  (
    .DIN(WX8616),
    .DIN_t(WX8616_t),
    .SDIN(n7717),
    .SDIN_t(n7717_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7718),
    .Q_t(n7718_t),
    .QN(n5242),
    .QN_t(n5242_t)
  );


  sdffs1
  \DFF_1290/Q_reg 
  (
    .DIN(WX8614),
    .DIN_t(WX8614_t),
    .SDIN(n7716),
    .SDIN_t(n7716_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7717),
    .Q_t(n7717_t),
    .QN(n5247),
    .QN_t(n5247_t)
  );


  sdffs1
  \DFF_1289/Q_reg 
  (
    .DIN(WX8612),
    .DIN_t(WX8612_t),
    .SDIN(n7715),
    .SDIN_t(n7715_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7716),
    .Q_t(n7716_t),
    .QN(n5252),
    .QN_t(n5252_t)
  );


  sdffs1
  \DFF_1288/Q_reg 
  (
    .DIN(WX8610),
    .DIN_t(WX8610_t),
    .SDIN(n7714),
    .SDIN_t(n7714_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7715),
    .Q_t(n7715_t),
    .QN(n5257),
    .QN_t(n5257_t)
  );


  sdffs1
  \DFF_1287/Q_reg 
  (
    .DIN(WX8608),
    .DIN_t(WX8608_t),
    .SDIN(n7713),
    .SDIN_t(n7713_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7714),
    .Q_t(n7714_t),
    .QN(n5262),
    .QN_t(n5262_t)
  );


  sdffs1
  \DFF_1286/Q_reg 
  (
    .DIN(WX8606),
    .DIN_t(WX8606_t),
    .SDIN(n7712),
    .SDIN_t(n7712_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7713),
    .Q_t(n7713_t),
    .QN(n5267),
    .QN_t(n5267_t)
  );


  sdffs1
  \DFF_1285/Q_reg 
  (
    .DIN(WX8604),
    .DIN_t(WX8604_t),
    .SDIN(n7711),
    .SDIN_t(n7711_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7712),
    .Q_t(n7712_t),
    .QN(n5272),
    .QN_t(n5272_t)
  );


  sdffs1
  \DFF_1284/Q_reg 
  (
    .DIN(WX8602),
    .DIN_t(WX8602_t),
    .SDIN(n7710),
    .SDIN_t(n7710_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7711),
    .Q_t(n7711_t),
    .QN(n5277),
    .QN_t(n5277_t)
  );


  sdffs1
  \DFF_1283/Q_reg 
  (
    .DIN(WX8600),
    .DIN_t(WX8600_t),
    .SDIN(n7709),
    .SDIN_t(n7709_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7710),
    .Q_t(n7710_t),
    .QN(n5282),
    .QN_t(n5282_t)
  );


  sdffs1
  \DFF_1282/Q_reg 
  (
    .DIN(WX8598),
    .DIN_t(WX8598_t),
    .SDIN(n7708),
    .SDIN_t(n7708_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7709),
    .Q_t(n7709_t),
    .QN(n5287),
    .QN_t(n5287_t)
  );


  sdffs1
  \DFF_1281/Q_reg 
  (
    .DIN(WX8596),
    .DIN_t(WX8596_t),
    .SDIN(n7707),
    .SDIN_t(n7707_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7708),
    .Q_t(n7708_t),
    .QN(n5292),
    .QN_t(n5292_t)
  );


  sdffs1
  \DFF_1280/Q_reg 
  (
    .DIN(WX8594),
    .DIN_t(WX8594_t),
    .SDIN(n7706),
    .SDIN_t(n7706_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7707),
    .Q_t(n7707_t),
    .QN(n5297),
    .QN_t(n5297_t)
  );


  sdffs1
  \DFF_1279/Q_reg 
  (
    .DIN(WX8592),
    .DIN_t(WX8592_t),
    .SDIN(n7705),
    .SDIN_t(n7705_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7706),
    .Q_t(n7706_t),
    .QN(n5157),
    .QN_t(n5157_t)
  );


  sdffs1
  \DFF_1278/Q_reg 
  (
    .DIN(WX8590),
    .DIN_t(WX8590_t),
    .SDIN(n7704),
    .SDIN_t(n7704_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7705),
    .Q_t(n7705_t),
    .QN(n5161),
    .QN_t(n5161_t)
  );


  sdffs1
  \DFF_1277/Q_reg 
  (
    .DIN(WX8588),
    .DIN_t(WX8588_t),
    .SDIN(n7703),
    .SDIN_t(n7703_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7704),
    .Q_t(n7704_t),
    .QN(n5165),
    .QN_t(n5165_t)
  );


  sdffs1
  \DFF_1276/Q_reg 
  (
    .DIN(WX8586),
    .DIN_t(WX8586_t),
    .SDIN(n7702),
    .SDIN_t(n7702_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7703),
    .Q_t(n7703_t),
    .QN(n5169),
    .QN_t(n5169_t)
  );


  sdffs1
  \DFF_1275/Q_reg 
  (
    .DIN(WX8584),
    .DIN_t(WX8584_t),
    .SDIN(n7701),
    .SDIN_t(n7701_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7702),
    .Q_t(n7702_t),
    .QN(n5173),
    .QN_t(n5173_t)
  );


  sdffs1
  \DFF_1274/Q_reg 
  (
    .DIN(WX8582),
    .DIN_t(WX8582_t),
    .SDIN(n7700),
    .SDIN_t(n7700_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7701),
    .Q_t(n7701_t),
    .QN(n5177),
    .QN_t(n5177_t)
  );


  sdffs1
  \DFF_1273/Q_reg 
  (
    .DIN(WX8580),
    .DIN_t(WX8580_t),
    .SDIN(n7699),
    .SDIN_t(n7699_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7700),
    .Q_t(n7700_t),
    .QN(n5181),
    .QN_t(n5181_t)
  );


  sdffs1
  \DFF_1272/Q_reg 
  (
    .DIN(WX8578),
    .DIN_t(WX8578_t),
    .SDIN(n7698),
    .SDIN_t(n7698_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7699),
    .Q_t(n7699_t),
    .QN(n5185),
    .QN_t(n5185_t)
  );


  sdffs1
  \DFF_1271/Q_reg 
  (
    .DIN(WX8576),
    .DIN_t(WX8576_t),
    .SDIN(n7697),
    .SDIN_t(n7697_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7698),
    .Q_t(n7698_t),
    .QN(n5189),
    .QN_t(n5189_t)
  );


  sdffs1
  \DFF_1270/Q_reg 
  (
    .DIN(WX8574),
    .DIN_t(WX8574_t),
    .SDIN(n7696),
    .SDIN_t(n7696_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7697),
    .Q_t(n7697_t),
    .QN(n5193),
    .QN_t(n5193_t)
  );


  sdffs1
  \DFF_1269/Q_reg 
  (
    .DIN(WX8572),
    .DIN_t(WX8572_t),
    .SDIN(n7695),
    .SDIN_t(n7695_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7696),
    .Q_t(n7696_t),
    .QN(n5197),
    .QN_t(n5197_t)
  );


  sdffs1
  \DFF_1268/Q_reg 
  (
    .DIN(WX8570),
    .DIN_t(WX8570_t),
    .SDIN(n7694),
    .SDIN_t(n7694_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7695),
    .Q_t(n7695_t),
    .QN(n5201),
    .QN_t(n5201_t)
  );


  sdffs1
  \DFF_1267/Q_reg 
  (
    .DIN(WX8568),
    .DIN_t(WX8568_t),
    .SDIN(n7693),
    .SDIN_t(n7693_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7694),
    .Q_t(n7694_t),
    .QN(n5205),
    .QN_t(n5205_t)
  );


  sdffs1
  \DFF_1266/Q_reg 
  (
    .DIN(WX8566),
    .DIN_t(WX8566_t),
    .SDIN(n7692),
    .SDIN_t(n7692_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7693),
    .Q_t(n7693_t),
    .QN(n5209),
    .QN_t(n5209_t)
  );


  sdffs1
  \DFF_1265/Q_reg 
  (
    .DIN(WX8564),
    .DIN_t(WX8564_t),
    .SDIN(n7691),
    .SDIN_t(n7691_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7692),
    .Q_t(n7692_t),
    .QN(n5213),
    .QN_t(n5213_t)
  );


  sdffs1
  \DFF_1264/Q_reg 
  (
    .DIN(WX8562),
    .DIN_t(WX8562_t),
    .SDIN(n7690),
    .SDIN_t(n7690_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7691),
    .Q_t(n7691_t),
    .QN(n5217),
    .QN_t(n5217_t)
  );


  sdffs1
  \DFF_1263/Q_reg 
  (
    .DIN(WX8560),
    .DIN_t(WX8560_t),
    .SDIN(n7689),
    .SDIN_t(n7689_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7690),
    .Q_t(n7690_t),
    .QN(n5221),
    .QN_t(n5221_t)
  );


  sdffs1
  \DFF_1262/Q_reg 
  (
    .DIN(WX8558),
    .DIN_t(WX8558_t),
    .SDIN(n7688),
    .SDIN_t(n7688_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7689),
    .Q_t(n7689_t),
    .QN(n5226),
    .QN_t(n5226_t)
  );


  sdffs1
  \DFF_1261/Q_reg 
  (
    .DIN(WX8556),
    .DIN_t(WX8556_t),
    .SDIN(n7687),
    .SDIN_t(n7687_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7688),
    .Q_t(n7688_t),
    .QN(n5231),
    .QN_t(n5231_t)
  );


  sdffs1
  \DFF_1260/Q_reg 
  (
    .DIN(WX8554),
    .DIN_t(WX8554_t),
    .SDIN(n7686),
    .SDIN_t(n7686_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7687),
    .Q_t(n7687_t),
    .QN(n5236),
    .QN_t(n5236_t)
  );


  sdffs1
  \DFF_1259/Q_reg 
  (
    .DIN(WX8552),
    .DIN_t(WX8552_t),
    .SDIN(n7685),
    .SDIN_t(n7685_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7686),
    .Q_t(n7686_t),
    .QN(n5241),
    .QN_t(n5241_t)
  );


  sdffs1
  \DFF_1258/Q_reg 
  (
    .DIN(WX8550),
    .DIN_t(WX8550_t),
    .SDIN(n7684),
    .SDIN_t(n7684_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7685),
    .Q_t(n7685_t),
    .QN(n5246),
    .QN_t(n5246_t)
  );


  sdffs1
  \DFF_1257/Q_reg 
  (
    .DIN(WX8548),
    .DIN_t(WX8548_t),
    .SDIN(n7683),
    .SDIN_t(n7683_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7684),
    .Q_t(n7684_t),
    .QN(n5251),
    .QN_t(n5251_t)
  );


  sdffs1
  \DFF_1256/Q_reg 
  (
    .DIN(WX8546),
    .DIN_t(WX8546_t),
    .SDIN(n7682),
    .SDIN_t(n7682_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7683),
    .Q_t(n7683_t),
    .QN(n5256),
    .QN_t(n5256_t)
  );


  sdffs1
  \DFF_1255/Q_reg 
  (
    .DIN(WX8544),
    .DIN_t(WX8544_t),
    .SDIN(n7681),
    .SDIN_t(n7681_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7682),
    .Q_t(n7682_t),
    .QN(n5261),
    .QN_t(n5261_t)
  );


  sdffs1
  \DFF_1254/Q_reg 
  (
    .DIN(WX8542),
    .DIN_t(WX8542_t),
    .SDIN(n7680),
    .SDIN_t(n7680_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7681),
    .Q_t(n7681_t),
    .QN(n5266),
    .QN_t(n5266_t)
  );


  sdffs1
  \DFF_1253/Q_reg 
  (
    .DIN(WX8540),
    .DIN_t(WX8540_t),
    .SDIN(n7679),
    .SDIN_t(n7679_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7680),
    .Q_t(n7680_t),
    .QN(n5271),
    .QN_t(n5271_t)
  );


  sdffs1
  \DFF_1252/Q_reg 
  (
    .DIN(WX8538),
    .DIN_t(WX8538_t),
    .SDIN(n7678),
    .SDIN_t(n7678_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7679),
    .Q_t(n7679_t),
    .QN(n5276),
    .QN_t(n5276_t)
  );


  sdffs1
  \DFF_1251/Q_reg 
  (
    .DIN(WX8536),
    .DIN_t(WX8536_t),
    .SDIN(n7677),
    .SDIN_t(n7677_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7678),
    .Q_t(n7678_t),
    .QN(n5281),
    .QN_t(n5281_t)
  );


  sdffs1
  \DFF_1250/Q_reg 
  (
    .DIN(WX8534),
    .DIN_t(WX8534_t),
    .SDIN(n7676),
    .SDIN_t(n7676_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7677),
    .Q_t(n7677_t),
    .QN(n5286),
    .QN_t(n5286_t)
  );


  sdffs1
  \DFF_1249/Q_reg 
  (
    .DIN(WX8532),
    .DIN_t(WX8532_t),
    .SDIN(n7675),
    .SDIN_t(n7675_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7676),
    .Q_t(n7676_t),
    .QN(n5291),
    .QN_t(n5291_t)
  );


  sdffs1
  \DFF_1248/Q_reg 
  (
    .DIN(WX8530),
    .DIN_t(WX8530_t),
    .SDIN(n7674),
    .SDIN_t(n7674_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7675),
    .Q_t(n7675_t),
    .QN(n5296),
    .QN_t(n5296_t)
  );


  sdffs1
  \DFF_1247/Q_reg 
  (
    .DIN(WX8528),
    .DIN_t(WX8528_t),
    .SDIN(n7673),
    .SDIN_t(n7673_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7674),
    .Q_t(n7674_t),
    .QN(n5156),
    .QN_t(n5156_t)
  );


  sdffs1
  \DFF_1246/Q_reg 
  (
    .DIN(WX8526),
    .DIN_t(WX8526_t),
    .SDIN(n7672),
    .SDIN_t(n7672_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7673),
    .Q_t(n7673_t),
    .QN(n5160),
    .QN_t(n5160_t)
  );


  sdffs1
  \DFF_1245/Q_reg 
  (
    .DIN(WX8524),
    .DIN_t(WX8524_t),
    .SDIN(n7671),
    .SDIN_t(n7671_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7672),
    .Q_t(n7672_t),
    .QN(n5164),
    .QN_t(n5164_t)
  );


  sdffs1
  \DFF_1244/Q_reg 
  (
    .DIN(WX8522),
    .DIN_t(WX8522_t),
    .SDIN(n7670),
    .SDIN_t(n7670_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7671),
    .Q_t(n7671_t),
    .QN(n5168),
    .QN_t(n5168_t)
  );


  sdffs1
  \DFF_1243/Q_reg 
  (
    .DIN(WX8520),
    .DIN_t(WX8520_t),
    .SDIN(n7669),
    .SDIN_t(n7669_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7670),
    .Q_t(n7670_t),
    .QN(n5172),
    .QN_t(n5172_t)
  );


  sdffs1
  \DFF_1242/Q_reg 
  (
    .DIN(WX8518),
    .DIN_t(WX8518_t),
    .SDIN(n7668),
    .SDIN_t(n7668_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7669),
    .Q_t(n7669_t),
    .QN(n5176),
    .QN_t(n5176_t)
  );


  sdffs1
  \DFF_1241/Q_reg 
  (
    .DIN(WX8516),
    .DIN_t(WX8516_t),
    .SDIN(n7667),
    .SDIN_t(n7667_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7668),
    .Q_t(n7668_t),
    .QN(n5180),
    .QN_t(n5180_t)
  );


  sdffs1
  \DFF_1240/Q_reg 
  (
    .DIN(WX8514),
    .DIN_t(WX8514_t),
    .SDIN(n7666),
    .SDIN_t(n7666_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7667),
    .Q_t(n7667_t),
    .QN(n5184),
    .QN_t(n5184_t)
  );


  sdffs1
  \DFF_1239/Q_reg 
  (
    .DIN(WX8512),
    .DIN_t(WX8512_t),
    .SDIN(n7665),
    .SDIN_t(n7665_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7666),
    .Q_t(n7666_t),
    .QN(n5188),
    .QN_t(n5188_t)
  );


  sdffs1
  \DFF_1238/Q_reg 
  (
    .DIN(WX8510),
    .DIN_t(WX8510_t),
    .SDIN(n7664),
    .SDIN_t(n7664_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7665),
    .Q_t(n7665_t),
    .QN(n5192),
    .QN_t(n5192_t)
  );


  sdffs1
  \DFF_1237/Q_reg 
  (
    .DIN(WX8508),
    .DIN_t(WX8508_t),
    .SDIN(n7663),
    .SDIN_t(n7663_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7664),
    .Q_t(n7664_t),
    .QN(n5196),
    .QN_t(n5196_t)
  );


  sdffs1
  \DFF_1236/Q_reg 
  (
    .DIN(WX8506),
    .DIN_t(WX8506_t),
    .SDIN(n7662),
    .SDIN_t(n7662_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7663),
    .Q_t(n7663_t),
    .QN(n5200),
    .QN_t(n5200_t)
  );


  sdffs1
  \DFF_1235/Q_reg 
  (
    .DIN(WX8504),
    .DIN_t(WX8504_t),
    .SDIN(n7661),
    .SDIN_t(n7661_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7662),
    .Q_t(n7662_t),
    .QN(n5204),
    .QN_t(n5204_t)
  );


  sdffs1
  \DFF_1234/Q_reg 
  (
    .DIN(WX8502),
    .DIN_t(WX8502_t),
    .SDIN(n7660),
    .SDIN_t(n7660_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7661),
    .Q_t(n7661_t),
    .QN(n5208),
    .QN_t(n5208_t)
  );


  sdffs1
  \DFF_1233/Q_reg 
  (
    .DIN(WX8500),
    .DIN_t(WX8500_t),
    .SDIN(n7659),
    .SDIN_t(n7659_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7660),
    .Q_t(n7660_t),
    .QN(n5212),
    .QN_t(n5212_t)
  );


  sdffs1
  \DFF_1232/Q_reg 
  (
    .DIN(WX8498),
    .DIN_t(WX8498_t),
    .SDIN(n5220),
    .SDIN_t(n5220_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7659),
    .Q_t(n7659_t),
    .QN(n5216),
    .QN_t(n5216_t)
  );


  sdffs1
  \DFF_1231/Q_reg 
  (
    .DIN(WX8496),
    .DIN_t(WX8496_t),
    .SDIN(n5225),
    .SDIN_t(n5225_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5220),
    .Q_t(n5220_t)
  );


  sdffs1
  \DFF_1230/Q_reg 
  (
    .DIN(WX8494),
    .DIN_t(WX8494_t),
    .SDIN(n5230),
    .SDIN_t(n5230_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5225),
    .Q_t(n5225_t)
  );


  sdffs1
  \DFF_1229/Q_reg 
  (
    .DIN(WX8492),
    .DIN_t(WX8492_t),
    .SDIN(n5235),
    .SDIN_t(n5235_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5230),
    .Q_t(n5230_t)
  );


  sdffs1
  \DFF_1228/Q_reg 
  (
    .DIN(WX8490),
    .DIN_t(WX8490_t),
    .SDIN(n5240),
    .SDIN_t(n5240_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5235),
    .Q_t(n5235_t)
  );


  sdffs1
  \DFF_1227/Q_reg 
  (
    .DIN(WX8488),
    .DIN_t(WX8488_t),
    .SDIN(n5245),
    .SDIN_t(n5245_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5240),
    .Q_t(n5240_t)
  );


  sdffs1
  \DFF_1226/Q_reg 
  (
    .DIN(WX8486),
    .DIN_t(WX8486_t),
    .SDIN(n5250),
    .SDIN_t(n5250_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5245),
    .Q_t(n5245_t)
  );


  sdffs1
  \DFF_1225/Q_reg 
  (
    .DIN(WX8484),
    .DIN_t(WX8484_t),
    .SDIN(n5255),
    .SDIN_t(n5255_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5250),
    .Q_t(n5250_t)
  );


  sdffs1
  \DFF_1224/Q_reg 
  (
    .DIN(WX8482),
    .DIN_t(WX8482_t),
    .SDIN(n5260),
    .SDIN_t(n5260_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5255),
    .Q_t(n5255_t)
  );


  sdffs1
  \DFF_1223/Q_reg 
  (
    .DIN(WX8480),
    .DIN_t(WX8480_t),
    .SDIN(n5265),
    .SDIN_t(n5265_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5260),
    .Q_t(n5260_t)
  );


  sdffs1
  \DFF_1222/Q_reg 
  (
    .DIN(WX8478),
    .DIN_t(WX8478_t),
    .SDIN(n5270),
    .SDIN_t(n5270_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5265),
    .Q_t(n5265_t)
  );


  sdffs1
  \DFF_1221/Q_reg 
  (
    .DIN(WX8476),
    .DIN_t(WX8476_t),
    .SDIN(n5275),
    .SDIN_t(n5275_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5270),
    .Q_t(n5270_t)
  );


  sdffs1
  \DFF_1220/Q_reg 
  (
    .DIN(WX8474),
    .DIN_t(WX8474_t),
    .SDIN(n5280),
    .SDIN_t(n5280_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5275),
    .Q_t(n5275_t)
  );


  sdffs1
  \DFF_1219/Q_reg 
  (
    .DIN(WX8472),
    .DIN_t(WX8472_t),
    .SDIN(n5285),
    .SDIN_t(n5285_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5280),
    .Q_t(n5280_t)
  );


  sdffs1
  \DFF_1218/Q_reg 
  (
    .DIN(WX8470),
    .DIN_t(WX8470_t),
    .SDIN(n5290),
    .SDIN_t(n5290_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5285),
    .Q_t(n5285_t)
  );


  sdffs1
  \DFF_1217/Q_reg 
  (
    .DIN(WX8468),
    .DIN_t(WX8468_t),
    .SDIN(n5295),
    .SDIN_t(n5295_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5290),
    .Q_t(n5290_t)
  );


  sdffs1
  \DFF_1216/Q_reg 
  (
    .DIN(WX8466),
    .DIN_t(WX8466_t),
    .SDIN(n5155),
    .SDIN_t(n5155_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5295),
    .Q_t(n5295_t)
  );


  sdffs1
  \DFF_1215/Q_reg 
  (
    .DIN(WX8464),
    .DIN_t(WX8464_t),
    .SDIN(n5159),
    .SDIN_t(n5159_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5155),
    .Q_t(n5155_t)
  );


  sdffs1
  \DFF_1214/Q_reg 
  (
    .DIN(WX8462),
    .DIN_t(WX8462_t),
    .SDIN(n5163),
    .SDIN_t(n5163_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5159),
    .Q_t(n5159_t)
  );


  sdffs1
  \DFF_1213/Q_reg 
  (
    .DIN(WX8460),
    .DIN_t(WX8460_t),
    .SDIN(n5167),
    .SDIN_t(n5167_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5163),
    .Q_t(n5163_t)
  );


  sdffs1
  \DFF_1212/Q_reg 
  (
    .DIN(WX8458),
    .DIN_t(WX8458_t),
    .SDIN(n5171),
    .SDIN_t(n5171_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5167),
    .Q_t(n5167_t)
  );


  sdffs1
  \DFF_1211/Q_reg 
  (
    .DIN(WX8456),
    .DIN_t(WX8456_t),
    .SDIN(n5175),
    .SDIN_t(n5175_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5171),
    .Q_t(n5171_t)
  );


  sdffs1
  \DFF_1210/Q_reg 
  (
    .DIN(WX8454),
    .DIN_t(WX8454_t),
    .SDIN(n5179),
    .SDIN_t(n5179_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5175),
    .Q_t(n5175_t)
  );


  sdffs1
  \DFF_1209/Q_reg 
  (
    .DIN(WX8452),
    .DIN_t(WX8452_t),
    .SDIN(n5183),
    .SDIN_t(n5183_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5179),
    .Q_t(n5179_t)
  );


  sdffs1
  \DFF_1208/Q_reg 
  (
    .DIN(WX8450),
    .DIN_t(WX8450_t),
    .SDIN(n5187),
    .SDIN_t(n5187_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5183),
    .Q_t(n5183_t)
  );


  sdffs1
  \DFF_1207/Q_reg 
  (
    .DIN(WX8448),
    .DIN_t(WX8448_t),
    .SDIN(n5191),
    .SDIN_t(n5191_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5187),
    .Q_t(n5187_t)
  );


  sdffs1
  \DFF_1206/Q_reg 
  (
    .DIN(WX8446),
    .DIN_t(WX8446_t),
    .SDIN(n5195),
    .SDIN_t(n5195_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5191),
    .Q_t(n5191_t)
  );


  sdffs1
  \DFF_1205/Q_reg 
  (
    .DIN(WX8444),
    .DIN_t(WX8444_t),
    .SDIN(n5199),
    .SDIN_t(n5199_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5195),
    .Q_t(n5195_t)
  );


  sdffs1
  \DFF_1204/Q_reg 
  (
    .DIN(WX8442),
    .DIN_t(WX8442_t),
    .SDIN(n5203),
    .SDIN_t(n5203_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5199),
    .Q_t(n5199_t)
  );


  sdffs1
  \DFF_1203/Q_reg 
  (
    .DIN(WX8440),
    .DIN_t(WX8440_t),
    .SDIN(n5207),
    .SDIN_t(n5207_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5203),
    .Q_t(n5203_t)
  );


  sdffs1
  \DFF_1202/Q_reg 
  (
    .DIN(WX8438),
    .DIN_t(WX8438_t),
    .SDIN(n5211),
    .SDIN_t(n5211_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5207),
    .Q_t(n5207_t)
  );


  sdffs1
  \DFF_1201/Q_reg 
  (
    .DIN(WX8436),
    .DIN_t(WX8436_t),
    .SDIN(n5215),
    .SDIN_t(n5215_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5211),
    .Q_t(n5211_t)
  );


  sdffs1
  \DFF_1200/Q_reg 
  (
    .DIN(WX8434),
    .DIN_t(WX8434_t),
    .SDIN(n7658),
    .SDIN_t(n7658_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5215),
    .Q_t(n5215_t)
  );


  sdffs1
  \DFF_1199/Q_reg 
  (
    .DIN(WX8432),
    .DIN_t(WX8432_t),
    .SDIN(n7657),
    .SDIN_t(n7657_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7658),
    .Q_t(n7658_t),
    .QN(n5219),
    .QN_t(n5219_t)
  );


  sdffs1
  \DFF_1198/Q_reg 
  (
    .DIN(WX8430),
    .DIN_t(WX8430_t),
    .SDIN(n7656),
    .SDIN_t(n7656_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7657),
    .Q_t(n7657_t),
    .QN(n5224),
    .QN_t(n5224_t)
  );


  sdffs1
  \DFF_1197/Q_reg 
  (
    .DIN(WX8428),
    .DIN_t(WX8428_t),
    .SDIN(n7655),
    .SDIN_t(n7655_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7656),
    .Q_t(n7656_t),
    .QN(n5229),
    .QN_t(n5229_t)
  );


  sdffs1
  \DFF_1196/Q_reg 
  (
    .DIN(WX8426),
    .DIN_t(WX8426_t),
    .SDIN(n7654),
    .SDIN_t(n7654_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7655),
    .Q_t(n7655_t),
    .QN(n5234),
    .QN_t(n5234_t)
  );


  sdffs1
  \DFF_1195/Q_reg 
  (
    .DIN(WX8424),
    .DIN_t(WX8424_t),
    .SDIN(n7653),
    .SDIN_t(n7653_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7654),
    .Q_t(n7654_t),
    .QN(n5239),
    .QN_t(n5239_t)
  );


  sdffs1
  \DFF_1194/Q_reg 
  (
    .DIN(WX8422),
    .DIN_t(WX8422_t),
    .SDIN(n7652),
    .SDIN_t(n7652_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7653),
    .Q_t(n7653_t),
    .QN(n5244),
    .QN_t(n5244_t)
  );


  sdffs1
  \DFF_1193/Q_reg 
  (
    .DIN(WX8420),
    .DIN_t(WX8420_t),
    .SDIN(n7651),
    .SDIN_t(n7651_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7652),
    .Q_t(n7652_t),
    .QN(n5249),
    .QN_t(n5249_t)
  );


  sdffs1
  \DFF_1192/Q_reg 
  (
    .DIN(WX8418),
    .DIN_t(WX8418_t),
    .SDIN(n7650),
    .SDIN_t(n7650_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7651),
    .Q_t(n7651_t),
    .QN(n5254),
    .QN_t(n5254_t)
  );


  sdffs1
  \DFF_1191/Q_reg 
  (
    .DIN(WX8416),
    .DIN_t(WX8416_t),
    .SDIN(n7649),
    .SDIN_t(n7649_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7650),
    .Q_t(n7650_t),
    .QN(n5259),
    .QN_t(n5259_t)
  );


  sdffs1
  \DFF_1190/Q_reg 
  (
    .DIN(WX8414),
    .DIN_t(WX8414_t),
    .SDIN(n7648),
    .SDIN_t(n7648_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7649),
    .Q_t(n7649_t),
    .QN(n5264),
    .QN_t(n5264_t)
  );


  sdffs1
  \DFF_1189/Q_reg 
  (
    .DIN(WX8412),
    .DIN_t(WX8412_t),
    .SDIN(n7647),
    .SDIN_t(n7647_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7648),
    .Q_t(n7648_t),
    .QN(n5269),
    .QN_t(n5269_t)
  );


  sdffs1
  \DFF_1188/Q_reg 
  (
    .DIN(WX8410),
    .DIN_t(WX8410_t),
    .SDIN(n7646),
    .SDIN_t(n7646_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7647),
    .Q_t(n7647_t),
    .QN(n5274),
    .QN_t(n5274_t)
  );


  sdffs1
  \DFF_1187/Q_reg 
  (
    .DIN(WX8408),
    .DIN_t(WX8408_t),
    .SDIN(n7645),
    .SDIN_t(n7645_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7646),
    .Q_t(n7646_t),
    .QN(n5279),
    .QN_t(n5279_t)
  );


  sdffs1
  \DFF_1186/Q_reg 
  (
    .DIN(WX8406),
    .DIN_t(WX8406_t),
    .SDIN(n7644),
    .SDIN_t(n7644_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7645),
    .Q_t(n7645_t),
    .QN(n5284),
    .QN_t(n5284_t)
  );


  sdffs1
  \DFF_1185/Q_reg 
  (
    .DIN(WX8404),
    .DIN_t(WX8404_t),
    .SDIN(n7643),
    .SDIN_t(n7643_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7644),
    .Q_t(n7644_t),
    .QN(n5289),
    .QN_t(n5289_t)
  );


  sdffs1
  \DFF_1184/Q_reg 
  (
    .DIN(WX8402),
    .DIN_t(WX8402_t),
    .SDIN(n7642),
    .SDIN_t(n7642_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7643),
    .Q_t(n7643_t),
    .QN(n5294),
    .QN_t(n5294_t)
  );


  sdffs1
  \DFF_1183/Q_reg 
  (
    .DIN(WX8304),
    .DIN_t(WX8304_t),
    .SDIN(n7641),
    .SDIN_t(n7641_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7642),
    .Q_t(n7642_t),
    .QN(n5124),
    .QN_t(n5124_t)
  );


  sdffs1
  \DFF_1182/Q_reg 
  (
    .DIN(WX8302),
    .DIN_t(WX8302_t),
    .SDIN(n7640),
    .SDIN_t(n7640_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7641),
    .Q_t(n7641_t),
    .QN(n5125),
    .QN_t(n5125_t)
  );


  sdffs1
  \DFF_1181/Q_reg 
  (
    .DIN(WX8300),
    .DIN_t(WX8300_t),
    .SDIN(n7639),
    .SDIN_t(n7639_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7640),
    .Q_t(n7640_t),
    .QN(n5126),
    .QN_t(n5126_t)
  );


  sdffs1
  \DFF_1180/Q_reg 
  (
    .DIN(WX8298),
    .DIN_t(WX8298_t),
    .SDIN(n7638),
    .SDIN_t(n7638_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7639),
    .Q_t(n7639_t),
    .QN(n5127),
    .QN_t(n5127_t)
  );


  sdffs1
  \DFF_1179/Q_reg 
  (
    .DIN(WX8296),
    .DIN_t(WX8296_t),
    .SDIN(n7637),
    .SDIN_t(n7637_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7638),
    .Q_t(n7638_t),
    .QN(n5128),
    .QN_t(n5128_t)
  );


  sdffs1
  \DFF_1178/Q_reg 
  (
    .DIN(WX8294),
    .DIN_t(WX8294_t),
    .SDIN(n7636),
    .SDIN_t(n7636_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7637),
    .Q_t(n7637_t),
    .QN(n5129),
    .QN_t(n5129_t)
  );


  sdffs1
  \DFF_1177/Q_reg 
  (
    .DIN(WX8292),
    .DIN_t(WX8292_t),
    .SDIN(n7635),
    .SDIN_t(n7635_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7636),
    .Q_t(n7636_t),
    .QN(n5130),
    .QN_t(n5130_t)
  );


  sdffs1
  \DFF_1176/Q_reg 
  (
    .DIN(WX8290),
    .DIN_t(WX8290_t),
    .SDIN(n7634),
    .SDIN_t(n7634_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7635),
    .Q_t(n7635_t),
    .QN(n5131),
    .QN_t(n5131_t)
  );


  sdffs1
  \DFF_1175/Q_reg 
  (
    .DIN(WX8288),
    .DIN_t(WX8288_t),
    .SDIN(n7633),
    .SDIN_t(n7633_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7634),
    .Q_t(n7634_t),
    .QN(n5132),
    .QN_t(n5132_t)
  );


  sdffs1
  \DFF_1174/Q_reg 
  (
    .DIN(WX8286),
    .DIN_t(WX8286_t),
    .SDIN(n7632),
    .SDIN_t(n7632_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7633),
    .Q_t(n7633_t),
    .QN(n5133),
    .QN_t(n5133_t)
  );


  sdffs1
  \DFF_1173/Q_reg 
  (
    .DIN(WX8284),
    .DIN_t(WX8284_t),
    .SDIN(n7631),
    .SDIN_t(n7631_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7632),
    .Q_t(n7632_t),
    .QN(n5134),
    .QN_t(n5134_t)
  );


  sdffs1
  \DFF_1172/Q_reg 
  (
    .DIN(WX8282),
    .DIN_t(WX8282_t),
    .SDIN(n7630),
    .SDIN_t(n7630_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7631),
    .Q_t(n7631_t),
    .QN(n5135),
    .QN_t(n5135_t)
  );


  sdffs1
  \DFF_1171/Q_reg 
  (
    .DIN(WX8280),
    .DIN_t(WX8280_t),
    .SDIN(n7629),
    .SDIN_t(n7629_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7630),
    .Q_t(n7630_t),
    .QN(n5136),
    .QN_t(n5136_t)
  );


  sdffs1
  \DFF_1170/Q_reg 
  (
    .DIN(WX8278),
    .DIN_t(WX8278_t),
    .SDIN(n7628),
    .SDIN_t(n7628_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7629),
    .Q_t(n7629_t),
    .QN(n5137),
    .QN_t(n5137_t)
  );


  sdffs1
  \DFF_1169/Q_reg 
  (
    .DIN(WX8276),
    .DIN_t(WX8276_t),
    .SDIN(n7627),
    .SDIN_t(n7627_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7628),
    .Q_t(n7628_t),
    .QN(n5138),
    .QN_t(n5138_t)
  );


  sdffs1
  \DFF_1168/Q_reg 
  (
    .DIN(WX8274),
    .DIN_t(WX8274_t),
    .SDIN(n7626),
    .SDIN_t(n7626_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7627),
    .Q_t(n7627_t),
    .QN(n5139),
    .QN_t(n5139_t)
  );


  sdffs1
  \DFF_1167/Q_reg 
  (
    .DIN(WX8272),
    .DIN_t(WX8272_t),
    .SDIN(n7625),
    .SDIN_t(n7625_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7626),
    .Q_t(n7626_t),
    .QN(n5140),
    .QN_t(n5140_t)
  );


  sdffs1
  \DFF_1166/Q_reg 
  (
    .DIN(WX8270),
    .DIN_t(WX8270_t),
    .SDIN(n7624),
    .SDIN_t(n7624_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7625),
    .Q_t(n7625_t),
    .QN(n5141),
    .QN_t(n5141_t)
  );


  sdffs1
  \DFF_1165/Q_reg 
  (
    .DIN(WX8268),
    .DIN_t(WX8268_t),
    .SDIN(n7623),
    .SDIN_t(n7623_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7624),
    .Q_t(n7624_t),
    .QN(n5142),
    .QN_t(n5142_t)
  );


  sdffs1
  \DFF_1164/Q_reg 
  (
    .DIN(WX8266),
    .DIN_t(WX8266_t),
    .SDIN(n7622),
    .SDIN_t(n7622_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7623),
    .Q_t(n7623_t),
    .QN(n5143),
    .QN_t(n5143_t)
  );


  sdffs1
  \DFF_1163/Q_reg 
  (
    .DIN(WX8264),
    .DIN_t(WX8264_t),
    .SDIN(n7621),
    .SDIN_t(n7621_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7622),
    .Q_t(n7622_t),
    .QN(n5144),
    .QN_t(n5144_t)
  );


  sdffs1
  \DFF_1162/Q_reg 
  (
    .DIN(WX8262),
    .DIN_t(WX8262_t),
    .SDIN(n7620),
    .SDIN_t(n7620_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7621),
    .Q_t(n7621_t),
    .QN(n5145),
    .QN_t(n5145_t)
  );


  sdffs1
  \DFF_1161/Q_reg 
  (
    .DIN(WX8260),
    .DIN_t(WX8260_t),
    .SDIN(n7619),
    .SDIN_t(n7619_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7620),
    .Q_t(n7620_t),
    .QN(n5146),
    .QN_t(n5146_t)
  );


  sdffs1
  \DFF_1160/Q_reg 
  (
    .DIN(WX8258),
    .DIN_t(WX8258_t),
    .SDIN(n7618),
    .SDIN_t(n7618_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7619),
    .Q_t(n7619_t),
    .QN(n5147),
    .QN_t(n5147_t)
  );


  sdffs1
  \DFF_1159/Q_reg 
  (
    .DIN(WX8256),
    .DIN_t(WX8256_t),
    .SDIN(n7617),
    .SDIN_t(n7617_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7618),
    .Q_t(n7618_t),
    .QN(n5148),
    .QN_t(n5148_t)
  );


  sdffs1
  \DFF_1158/Q_reg 
  (
    .DIN(WX8254),
    .DIN_t(WX8254_t),
    .SDIN(n7616),
    .SDIN_t(n7616_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7617),
    .Q_t(n7617_t),
    .QN(n5149),
    .QN_t(n5149_t)
  );


  sdffs1
  \DFF_1157/Q_reg 
  (
    .DIN(WX8252),
    .DIN_t(WX8252_t),
    .SDIN(n7615),
    .SDIN_t(n7615_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7616),
    .Q_t(n7616_t),
    .QN(n5150),
    .QN_t(n5150_t)
  );


  sdffs1
  \DFF_1156/Q_reg 
  (
    .DIN(WX8250),
    .DIN_t(WX8250_t),
    .SDIN(n7614),
    .SDIN_t(n7614_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7615),
    .Q_t(n7615_t),
    .QN(n5151),
    .QN_t(n5151_t)
  );


  sdffs1
  \DFF_1155/Q_reg 
  (
    .DIN(WX8248),
    .DIN_t(WX8248_t),
    .SDIN(n7613),
    .SDIN_t(n7613_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7614),
    .Q_t(n7614_t),
    .QN(n5152),
    .QN_t(n5152_t)
  );


  sdffs1
  \DFF_1154/Q_reg 
  (
    .DIN(WX8246),
    .DIN_t(WX8246_t),
    .SDIN(n7612),
    .SDIN_t(n7612_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7613),
    .Q_t(n7613_t),
    .QN(n5153),
    .QN_t(n5153_t)
  );


  sdffs1
  \DFF_1153/Q_reg 
  (
    .DIN(WX8244),
    .DIN_t(WX8244_t),
    .SDIN(n7611),
    .SDIN_t(n7611_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7612),
    .Q_t(n7612_t),
    .QN(n5154),
    .QN_t(n5154_t)
  );


  sdffs1
  \DFF_1152/Q_reg 
  (
    .DIN(WX8242),
    .DIN_t(WX8242_t),
    .SDIN(CRC_OUT_4_31),
    .SDIN_t(CRC_OUT_4_31_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7611),
    .Q_t(n7611_t),
    .QN(n5123),
    .QN_t(n5123_t)
  );


  sdffs1
  \DFF_1151/Q_reg 
  (
    .DIN(WX7791),
    .DIN_t(WX7791_t),
    .SDIN(CRC_OUT_4_30),
    .SDIN_t(CRC_OUT_4_30_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_31),
    .Q_t(CRC_OUT_4_31_t),
    .QN(n5298),
    .QN_t(n5298_t)
  );


  sdffs1
  \DFF_1150/Q_reg 
  (
    .DIN(WX7789),
    .DIN_t(WX7789_t),
    .SDIN(CRC_OUT_4_29),
    .SDIN_t(CRC_OUT_4_29_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_30),
    .Q_t(CRC_OUT_4_30_t),
    .QN(n5293),
    .QN_t(n5293_t)
  );


  sdffs1
  \DFF_1149/Q_reg 
  (
    .DIN(WX7787),
    .DIN_t(WX7787_t),
    .SDIN(CRC_OUT_4_28),
    .SDIN_t(CRC_OUT_4_28_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_29),
    .Q_t(CRC_OUT_4_29_t),
    .QN(n5288),
    .QN_t(n5288_t)
  );


  sdffs1
  \DFF_1148/Q_reg 
  (
    .DIN(WX7785),
    .DIN_t(WX7785_t),
    .SDIN(CRC_OUT_4_27),
    .SDIN_t(CRC_OUT_4_27_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_28),
    .Q_t(CRC_OUT_4_28_t),
    .QN(n5283),
    .QN_t(n5283_t)
  );


  sdffs1
  \DFF_1147/Q_reg 
  (
    .DIN(WX7783),
    .DIN_t(WX7783_t),
    .SDIN(CRC_OUT_4_26),
    .SDIN_t(CRC_OUT_4_26_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_27),
    .Q_t(CRC_OUT_4_27_t),
    .QN(n5278),
    .QN_t(n5278_t)
  );


  sdffs1
  \DFF_1146/Q_reg 
  (
    .DIN(WX7781),
    .DIN_t(WX7781_t),
    .SDIN(CRC_OUT_4_25),
    .SDIN_t(CRC_OUT_4_25_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_26),
    .Q_t(CRC_OUT_4_26_t),
    .QN(n5273),
    .QN_t(n5273_t)
  );


  sdffs1
  \DFF_1145/Q_reg 
  (
    .DIN(WX7779),
    .DIN_t(WX7779_t),
    .SDIN(CRC_OUT_4_24),
    .SDIN_t(CRC_OUT_4_24_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_25),
    .Q_t(CRC_OUT_4_25_t),
    .QN(n5268),
    .QN_t(n5268_t)
  );


  sdffs1
  \DFF_1144/Q_reg 
  (
    .DIN(WX7777),
    .DIN_t(WX7777_t),
    .SDIN(CRC_OUT_4_23),
    .SDIN_t(CRC_OUT_4_23_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_24),
    .Q_t(CRC_OUT_4_24_t),
    .QN(n5263),
    .QN_t(n5263_t)
  );


  sdffs1
  \DFF_1143/Q_reg 
  (
    .DIN(WX7775),
    .DIN_t(WX7775_t),
    .SDIN(CRC_OUT_4_22),
    .SDIN_t(CRC_OUT_4_22_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_23),
    .Q_t(CRC_OUT_4_23_t),
    .QN(n5258),
    .QN_t(n5258_t)
  );


  sdffs1
  \DFF_1142/Q_reg 
  (
    .DIN(WX7773),
    .DIN_t(WX7773_t),
    .SDIN(CRC_OUT_4_21),
    .SDIN_t(CRC_OUT_4_21_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_22),
    .Q_t(CRC_OUT_4_22_t),
    .QN(n5253),
    .QN_t(n5253_t)
  );


  sdffs1
  \DFF_1141/Q_reg 
  (
    .DIN(WX7771),
    .DIN_t(WX7771_t),
    .SDIN(CRC_OUT_4_20),
    .SDIN_t(CRC_OUT_4_20_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_21),
    .Q_t(CRC_OUT_4_21_t),
    .QN(n5248),
    .QN_t(n5248_t)
  );


  sdffs1
  \DFF_1140/Q_reg 
  (
    .DIN(WX7769),
    .DIN_t(WX7769_t),
    .SDIN(CRC_OUT_4_19),
    .SDIN_t(CRC_OUT_4_19_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_20),
    .Q_t(CRC_OUT_4_20_t),
    .QN(n5243),
    .QN_t(n5243_t)
  );


  sdffs1
  \DFF_1139/Q_reg 
  (
    .DIN(WX7767),
    .DIN_t(WX7767_t),
    .SDIN(CRC_OUT_4_18),
    .SDIN_t(CRC_OUT_4_18_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_19),
    .Q_t(CRC_OUT_4_19_t),
    .QN(n5238),
    .QN_t(n5238_t)
  );


  sdffs1
  \DFF_1138/Q_reg 
  (
    .DIN(WX7765),
    .DIN_t(WX7765_t),
    .SDIN(CRC_OUT_4_17),
    .SDIN_t(CRC_OUT_4_17_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_18),
    .Q_t(CRC_OUT_4_18_t),
    .QN(n5233),
    .QN_t(n5233_t)
  );


  sdffs1
  \DFF_1137/Q_reg 
  (
    .DIN(WX7763),
    .DIN_t(WX7763_t),
    .SDIN(CRC_OUT_4_16),
    .SDIN_t(CRC_OUT_4_16_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_17),
    .Q_t(CRC_OUT_4_17_t),
    .QN(n5228),
    .QN_t(n5228_t)
  );


  sdffs1
  \DFF_1136/Q_reg 
  (
    .DIN(WX7761),
    .DIN_t(WX7761_t),
    .SDIN(CRC_OUT_4_15),
    .SDIN_t(CRC_OUT_4_15_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_16),
    .Q_t(CRC_OUT_4_16_t),
    .QN(n5223),
    .QN_t(n5223_t)
  );


  sdffs1
  \DFF_1135/Q_reg 
  (
    .DIN(WX7759),
    .DIN_t(WX7759_t),
    .SDIN(CRC_OUT_4_14),
    .SDIN_t(CRC_OUT_4_14_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_15),
    .Q_t(CRC_OUT_4_15_t),
    .QN(n5218),
    .QN_t(n5218_t)
  );


  sdffs1
  \DFF_1134/Q_reg 
  (
    .DIN(WX7757),
    .DIN_t(WX7757_t),
    .SDIN(CRC_OUT_4_13),
    .SDIN_t(CRC_OUT_4_13_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_14),
    .Q_t(CRC_OUT_4_14_t),
    .QN(n5214),
    .QN_t(n5214_t)
  );


  sdffs1
  \DFF_1133/Q_reg 
  (
    .DIN(WX7755),
    .DIN_t(WX7755_t),
    .SDIN(CRC_OUT_4_12),
    .SDIN_t(CRC_OUT_4_12_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_13),
    .Q_t(CRC_OUT_4_13_t),
    .QN(n5210),
    .QN_t(n5210_t)
  );


  sdffs1
  \DFF_1132/Q_reg 
  (
    .DIN(WX7753),
    .DIN_t(WX7753_t),
    .SDIN(CRC_OUT_4_11),
    .SDIN_t(CRC_OUT_4_11_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_12),
    .Q_t(CRC_OUT_4_12_t),
    .QN(n5206),
    .QN_t(n5206_t)
  );


  sdffs1
  \DFF_1131/Q_reg 
  (
    .DIN(WX7751),
    .DIN_t(WX7751_t),
    .SDIN(CRC_OUT_4_10),
    .SDIN_t(CRC_OUT_4_10_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_11),
    .Q_t(CRC_OUT_4_11_t),
    .QN(n5202),
    .QN_t(n5202_t)
  );


  sdffs1
  \DFF_1130/Q_reg 
  (
    .DIN(WX7749),
    .DIN_t(WX7749_t),
    .SDIN(CRC_OUT_4_9),
    .SDIN_t(CRC_OUT_4_9_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_10),
    .Q_t(CRC_OUT_4_10_t),
    .QN(n5198),
    .QN_t(n5198_t)
  );


  sdffs1
  \DFF_1129/Q_reg 
  (
    .DIN(WX7747),
    .DIN_t(WX7747_t),
    .SDIN(CRC_OUT_4_8),
    .SDIN_t(CRC_OUT_4_8_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_9),
    .Q_t(CRC_OUT_4_9_t),
    .QN(n5194),
    .QN_t(n5194_t)
  );


  sdffs1
  \DFF_1128/Q_reg 
  (
    .DIN(WX7745),
    .DIN_t(WX7745_t),
    .SDIN(CRC_OUT_4_7),
    .SDIN_t(CRC_OUT_4_7_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_8),
    .Q_t(CRC_OUT_4_8_t),
    .QN(n5190),
    .QN_t(n5190_t)
  );


  sdffs1
  \DFF_1127/Q_reg 
  (
    .DIN(WX7743),
    .DIN_t(WX7743_t),
    .SDIN(CRC_OUT_4_6),
    .SDIN_t(CRC_OUT_4_6_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_7),
    .Q_t(CRC_OUT_4_7_t),
    .QN(n5186),
    .QN_t(n5186_t)
  );


  sdffs1
  \DFF_1126/Q_reg 
  (
    .DIN(WX7741),
    .DIN_t(WX7741_t),
    .SDIN(CRC_OUT_4_5),
    .SDIN_t(CRC_OUT_4_5_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_6),
    .Q_t(CRC_OUT_4_6_t),
    .QN(n5182),
    .QN_t(n5182_t)
  );


  sdffs1
  \DFF_1125/Q_reg 
  (
    .DIN(WX7739),
    .DIN_t(WX7739_t),
    .SDIN(CRC_OUT_4_4),
    .SDIN_t(CRC_OUT_4_4_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_5),
    .Q_t(CRC_OUT_4_5_t),
    .QN(n5178),
    .QN_t(n5178_t)
  );


  sdffs1
  \DFF_1124/Q_reg 
  (
    .DIN(WX7737),
    .DIN_t(WX7737_t),
    .SDIN(CRC_OUT_4_3),
    .SDIN_t(CRC_OUT_4_3_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_4),
    .Q_t(CRC_OUT_4_4_t),
    .QN(n5174),
    .QN_t(n5174_t)
  );


  sdffs1
  \DFF_1123/Q_reg 
  (
    .DIN(WX7735),
    .DIN_t(WX7735_t),
    .SDIN(CRC_OUT_4_2),
    .SDIN_t(CRC_OUT_4_2_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_3),
    .Q_t(CRC_OUT_4_3_t),
    .QN(n5170),
    .QN_t(n5170_t)
  );


  sdffs1
  \DFF_1122/Q_reg 
  (
    .DIN(WX7733),
    .DIN_t(WX7733_t),
    .SDIN(CRC_OUT_4_1),
    .SDIN_t(CRC_OUT_4_1_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_2),
    .Q_t(CRC_OUT_4_2_t),
    .QN(n5166),
    .QN_t(n5166_t)
  );


  sdffs1
  \DFF_1121/Q_reg 
  (
    .DIN(WX7731),
    .DIN_t(WX7731_t),
    .SDIN(CRC_OUT_4_0),
    .SDIN_t(CRC_OUT_4_0_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_1),
    .Q_t(CRC_OUT_4_1_t),
    .QN(n5162),
    .QN_t(n5162_t)
  );


  sdffs1
  \DFF_1120/Q_reg 
  (
    .DIN(WX7729),
    .DIN_t(WX7729_t),
    .SDIN(n7610),
    .SDIN_t(n7610_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_4_0),
    .Q_t(CRC_OUT_4_0_t),
    .QN(n5158),
    .QN_t(n5158_t)
  );


  sdffs1
  \DFF_1119/Q_reg 
  (
    .DIN(WX7363),
    .DIN_t(WX7363_t),
    .SDIN(n7609),
    .SDIN_t(n7609_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7610),
    .Q_t(n7610_t),
    .QN(n3237),
    .QN_t(n3237_t)
  );


  sdffs1
  \DFF_1118/Q_reg 
  (
    .DIN(WX7361),
    .DIN_t(WX7361_t),
    .SDIN(n7608),
    .SDIN_t(n7608_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7609),
    .Q_t(n7609_t),
    .QN(n3238),
    .QN_t(n3238_t)
  );


  sdffs1
  \DFF_1117/Q_reg 
  (
    .DIN(WX7359),
    .DIN_t(WX7359_t),
    .SDIN(n7607),
    .SDIN_t(n7607_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7608),
    .Q_t(n7608_t),
    .QN(n3239),
    .QN_t(n3239_t)
  );


  sdffs1
  \DFF_1116/Q_reg 
  (
    .DIN(WX7357),
    .DIN_t(WX7357_t),
    .SDIN(n7606),
    .SDIN_t(n7606_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7607),
    .Q_t(n7607_t),
    .QN(n3240),
    .QN_t(n3240_t)
  );


  sdffs1
  \DFF_1115/Q_reg 
  (
    .DIN(WX7355),
    .DIN_t(WX7355_t),
    .SDIN(n7605),
    .SDIN_t(n7605_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7606),
    .Q_t(n7606_t),
    .QN(n3241),
    .QN_t(n3241_t)
  );


  sdffs1
  \DFF_1114/Q_reg 
  (
    .DIN(WX7353),
    .DIN_t(WX7353_t),
    .SDIN(n7604),
    .SDIN_t(n7604_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7605),
    .Q_t(n7605_t),
    .QN(n3242),
    .QN_t(n3242_t)
  );


  sdffs1
  \DFF_1113/Q_reg 
  (
    .DIN(WX7351),
    .DIN_t(WX7351_t),
    .SDIN(n7603),
    .SDIN_t(n7603_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7604),
    .Q_t(n7604_t),
    .QN(n3243),
    .QN_t(n3243_t)
  );


  sdffs1
  \DFF_1112/Q_reg 
  (
    .DIN(WX7349),
    .DIN_t(WX7349_t),
    .SDIN(n7602),
    .SDIN_t(n7602_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7603),
    .Q_t(n7603_t),
    .QN(n3244),
    .QN_t(n3244_t)
  );


  sdffs1
  \DFF_1111/Q_reg 
  (
    .DIN(WX7347),
    .DIN_t(WX7347_t),
    .SDIN(n7601),
    .SDIN_t(n7601_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7602),
    .Q_t(n7602_t),
    .QN(n3245),
    .QN_t(n3245_t)
  );


  sdffs1
  \DFF_1110/Q_reg 
  (
    .DIN(WX7345),
    .DIN_t(WX7345_t),
    .SDIN(n7600),
    .SDIN_t(n7600_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7601),
    .Q_t(n7601_t),
    .QN(n3246),
    .QN_t(n3246_t)
  );


  sdffs1
  \DFF_1109/Q_reg 
  (
    .DIN(WX7343),
    .DIN_t(WX7343_t),
    .SDIN(n7599),
    .SDIN_t(n7599_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7600),
    .Q_t(n7600_t),
    .QN(n3247),
    .QN_t(n3247_t)
  );


  sdffs1
  \DFF_1108/Q_reg 
  (
    .DIN(WX7341),
    .DIN_t(WX7341_t),
    .SDIN(n7598),
    .SDIN_t(n7598_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7599),
    .Q_t(n7599_t),
    .QN(n3248),
    .QN_t(n3248_t)
  );


  sdffs1
  \DFF_1107/Q_reg 
  (
    .DIN(WX7339),
    .DIN_t(WX7339_t),
    .SDIN(n7597),
    .SDIN_t(n7597_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7598),
    .Q_t(n7598_t),
    .QN(n3249),
    .QN_t(n3249_t)
  );


  sdffs1
  \DFF_1106/Q_reg 
  (
    .DIN(WX7337),
    .DIN_t(WX7337_t),
    .SDIN(n7596),
    .SDIN_t(n7596_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7597),
    .Q_t(n7597_t),
    .QN(n3250),
    .QN_t(n3250_t)
  );


  sdffs1
  \DFF_1105/Q_reg 
  (
    .DIN(WX7335),
    .DIN_t(WX7335_t),
    .SDIN(n7595),
    .SDIN_t(n7595_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7596),
    .Q_t(n7596_t),
    .QN(n3251),
    .QN_t(n3251_t)
  );


  sdffs1
  \DFF_1104/Q_reg 
  (
    .DIN(WX7333),
    .DIN_t(WX7333_t),
    .SDIN(n7594),
    .SDIN_t(n7594_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7595),
    .Q_t(n7595_t),
    .QN(n3252),
    .QN_t(n3252_t)
  );


  sdffs1
  \DFF_1103/Q_reg 
  (
    .DIN(WX7331),
    .DIN_t(WX7331_t),
    .SDIN(n7593),
    .SDIN_t(n7593_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7594),
    .Q_t(n7594_t),
    .QN(n5398),
    .QN_t(n5398_t)
  );


  sdffs1
  \DFF_1102/Q_reg 
  (
    .DIN(WX7329),
    .DIN_t(WX7329_t),
    .SDIN(n7592),
    .SDIN_t(n7592_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7593),
    .Q_t(n7593_t),
    .QN(n5403),
    .QN_t(n5403_t)
  );


  sdffs1
  \DFF_1101/Q_reg 
  (
    .DIN(WX7327),
    .DIN_t(WX7327_t),
    .SDIN(n7591),
    .SDIN_t(n7591_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7592),
    .Q_t(n7592_t),
    .QN(n5408),
    .QN_t(n5408_t)
  );


  sdffs1
  \DFF_1100/Q_reg 
  (
    .DIN(WX7325),
    .DIN_t(WX7325_t),
    .SDIN(n7590),
    .SDIN_t(n7590_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7591),
    .Q_t(n7591_t),
    .QN(n5413),
    .QN_t(n5413_t)
  );


  sdffs1
  \DFF_1099/Q_reg 
  (
    .DIN(WX7323),
    .DIN_t(WX7323_t),
    .SDIN(n7589),
    .SDIN_t(n7589_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7590),
    .Q_t(n7590_t),
    .QN(n5418),
    .QN_t(n5418_t)
  );


  sdffs1
  \DFF_1098/Q_reg 
  (
    .DIN(WX7321),
    .DIN_t(WX7321_t),
    .SDIN(n7588),
    .SDIN_t(n7588_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7589),
    .Q_t(n7589_t),
    .QN(n5423),
    .QN_t(n5423_t)
  );


  sdffs1
  \DFF_1097/Q_reg 
  (
    .DIN(WX7319),
    .DIN_t(WX7319_t),
    .SDIN(n7587),
    .SDIN_t(n7587_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7588),
    .Q_t(n7588_t),
    .QN(n5428),
    .QN_t(n5428_t)
  );


  sdffs1
  \DFF_1096/Q_reg 
  (
    .DIN(WX7317),
    .DIN_t(WX7317_t),
    .SDIN(n7586),
    .SDIN_t(n7586_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7587),
    .Q_t(n7587_t),
    .QN(n5433),
    .QN_t(n5433_t)
  );


  sdffs1
  \DFF_1095/Q_reg 
  (
    .DIN(WX7315),
    .DIN_t(WX7315_t),
    .SDIN(n7585),
    .SDIN_t(n7585_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7586),
    .Q_t(n7586_t),
    .QN(n5438),
    .QN_t(n5438_t)
  );


  sdffs1
  \DFF_1094/Q_reg 
  (
    .DIN(WX7313),
    .DIN_t(WX7313_t),
    .SDIN(n7584),
    .SDIN_t(n7584_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7585),
    .Q_t(n7585_t),
    .QN(n5443),
    .QN_t(n5443_t)
  );


  sdffs1
  \DFF_1093/Q_reg 
  (
    .DIN(WX7311),
    .DIN_t(WX7311_t),
    .SDIN(n7583),
    .SDIN_t(n7583_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7584),
    .Q_t(n7584_t),
    .QN(n5448),
    .QN_t(n5448_t)
  );


  sdffs1
  \DFF_1092/Q_reg 
  (
    .DIN(WX7309),
    .DIN_t(WX7309_t),
    .SDIN(n7582),
    .SDIN_t(n7582_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7583),
    .Q_t(n7583_t),
    .QN(n5453),
    .QN_t(n5453_t)
  );


  sdffs1
  \DFF_1091/Q_reg 
  (
    .DIN(WX7307),
    .DIN_t(WX7307_t),
    .SDIN(n7581),
    .SDIN_t(n7581_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7582),
    .Q_t(n7582_t),
    .QN(n5458),
    .QN_t(n5458_t)
  );


  sdffs1
  \DFF_1090/Q_reg 
  (
    .DIN(WX7305),
    .DIN_t(WX7305_t),
    .SDIN(n7580),
    .SDIN_t(n7580_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7581),
    .Q_t(n7581_t),
    .QN(n5463),
    .QN_t(n5463_t)
  );


  sdffs1
  \DFF_1089/Q_reg 
  (
    .DIN(WX7303),
    .DIN_t(WX7303_t),
    .SDIN(n7579),
    .SDIN_t(n7579_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7580),
    .Q_t(n7580_t),
    .QN(n5468),
    .QN_t(n5468_t)
  );


  sdffs1
  \DFF_1088/Q_reg 
  (
    .DIN(WX7301),
    .DIN_t(WX7301_t),
    .SDIN(n7578),
    .SDIN_t(n7578_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7579),
    .Q_t(n7579_t),
    .QN(n5473),
    .QN_t(n5473_t)
  );


  sdffs1
  \DFF_1087/Q_reg 
  (
    .DIN(WX7299),
    .DIN_t(WX7299_t),
    .SDIN(n7577),
    .SDIN_t(n7577_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7578),
    .Q_t(n7578_t),
    .QN(n5333),
    .QN_t(n5333_t)
  );


  sdffs1
  \DFF_1086/Q_reg 
  (
    .DIN(WX7297),
    .DIN_t(WX7297_t),
    .SDIN(n7576),
    .SDIN_t(n7576_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7577),
    .Q_t(n7577_t),
    .QN(n5337),
    .QN_t(n5337_t)
  );


  sdffs1
  \DFF_1085/Q_reg 
  (
    .DIN(WX7295),
    .DIN_t(WX7295_t),
    .SDIN(n7575),
    .SDIN_t(n7575_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7576),
    .Q_t(n7576_t),
    .QN(n5341),
    .QN_t(n5341_t)
  );


  sdffs1
  \DFF_1084/Q_reg 
  (
    .DIN(WX7293),
    .DIN_t(WX7293_t),
    .SDIN(n7574),
    .SDIN_t(n7574_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7575),
    .Q_t(n7575_t),
    .QN(n5345),
    .QN_t(n5345_t)
  );


  sdffs1
  \DFF_1083/Q_reg 
  (
    .DIN(WX7291),
    .DIN_t(WX7291_t),
    .SDIN(n7573),
    .SDIN_t(n7573_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7574),
    .Q_t(n7574_t),
    .QN(n5349),
    .QN_t(n5349_t)
  );


  sdffs1
  \DFF_1082/Q_reg 
  (
    .DIN(WX7289),
    .DIN_t(WX7289_t),
    .SDIN(n7572),
    .SDIN_t(n7572_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7573),
    .Q_t(n7573_t),
    .QN(n5353),
    .QN_t(n5353_t)
  );


  sdffs1
  \DFF_1081/Q_reg 
  (
    .DIN(WX7287),
    .DIN_t(WX7287_t),
    .SDIN(n7571),
    .SDIN_t(n7571_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7572),
    .Q_t(n7572_t),
    .QN(n5357),
    .QN_t(n5357_t)
  );


  sdffs1
  \DFF_1080/Q_reg 
  (
    .DIN(WX7285),
    .DIN_t(WX7285_t),
    .SDIN(n7570),
    .SDIN_t(n7570_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7571),
    .Q_t(n7571_t),
    .QN(n5361),
    .QN_t(n5361_t)
  );


  sdffs1
  \DFF_1079/Q_reg 
  (
    .DIN(WX7283),
    .DIN_t(WX7283_t),
    .SDIN(n7569),
    .SDIN_t(n7569_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7570),
    .Q_t(n7570_t),
    .QN(n5365),
    .QN_t(n5365_t)
  );


  sdffs1
  \DFF_1078/Q_reg 
  (
    .DIN(WX7281),
    .DIN_t(WX7281_t),
    .SDIN(n7568),
    .SDIN_t(n7568_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7569),
    .Q_t(n7569_t),
    .QN(n5369),
    .QN_t(n5369_t)
  );


  sdffs1
  \DFF_1077/Q_reg 
  (
    .DIN(WX7279),
    .DIN_t(WX7279_t),
    .SDIN(n7567),
    .SDIN_t(n7567_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7568),
    .Q_t(n7568_t),
    .QN(n5373),
    .QN_t(n5373_t)
  );


  sdffs1
  \DFF_1076/Q_reg 
  (
    .DIN(WX7277),
    .DIN_t(WX7277_t),
    .SDIN(n7566),
    .SDIN_t(n7566_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7567),
    .Q_t(n7567_t),
    .QN(n5377),
    .QN_t(n5377_t)
  );


  sdffs1
  \DFF_1075/Q_reg 
  (
    .DIN(WX7275),
    .DIN_t(WX7275_t),
    .SDIN(n7565),
    .SDIN_t(n7565_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7566),
    .Q_t(n7566_t),
    .QN(n5381),
    .QN_t(n5381_t)
  );


  sdffs1
  \DFF_1074/Q_reg 
  (
    .DIN(WX7273),
    .DIN_t(WX7273_t),
    .SDIN(n7564),
    .SDIN_t(n7564_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7565),
    .Q_t(n7565_t),
    .QN(n5385),
    .QN_t(n5385_t)
  );


  sdffs1
  \DFF_1073/Q_reg 
  (
    .DIN(WX7271),
    .DIN_t(WX7271_t),
    .SDIN(n7563),
    .SDIN_t(n7563_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7564),
    .Q_t(n7564_t),
    .QN(n5389),
    .QN_t(n5389_t)
  );


  sdffs1
  \DFF_1072/Q_reg 
  (
    .DIN(WX7269),
    .DIN_t(WX7269_t),
    .SDIN(n7562),
    .SDIN_t(n7562_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7563),
    .Q_t(n7563_t),
    .QN(n5393),
    .QN_t(n5393_t)
  );


  sdffs1
  \DFF_1071/Q_reg 
  (
    .DIN(WX7267),
    .DIN_t(WX7267_t),
    .SDIN(n7561),
    .SDIN_t(n7561_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7562),
    .Q_t(n7562_t),
    .QN(n5397),
    .QN_t(n5397_t)
  );


  sdffs1
  \DFF_1070/Q_reg 
  (
    .DIN(WX7265),
    .DIN_t(WX7265_t),
    .SDIN(n7560),
    .SDIN_t(n7560_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7561),
    .Q_t(n7561_t),
    .QN(n5402),
    .QN_t(n5402_t)
  );


  sdffs1
  \DFF_1069/Q_reg 
  (
    .DIN(WX7263),
    .DIN_t(WX7263_t),
    .SDIN(n7559),
    .SDIN_t(n7559_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7560),
    .Q_t(n7560_t),
    .QN(n5407),
    .QN_t(n5407_t)
  );


  sdffs1
  \DFF_1068/Q_reg 
  (
    .DIN(WX7261),
    .DIN_t(WX7261_t),
    .SDIN(n7558),
    .SDIN_t(n7558_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7559),
    .Q_t(n7559_t),
    .QN(n5412),
    .QN_t(n5412_t)
  );


  sdffs1
  \DFF_1067/Q_reg 
  (
    .DIN(WX7259),
    .DIN_t(WX7259_t),
    .SDIN(n7557),
    .SDIN_t(n7557_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7558),
    .Q_t(n7558_t),
    .QN(n5417),
    .QN_t(n5417_t)
  );


  sdffs1
  \DFF_1066/Q_reg 
  (
    .DIN(WX7257),
    .DIN_t(WX7257_t),
    .SDIN(n7556),
    .SDIN_t(n7556_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7557),
    .Q_t(n7557_t),
    .QN(n5422),
    .QN_t(n5422_t)
  );


  sdffs1
  \DFF_1065/Q_reg 
  (
    .DIN(WX7255),
    .DIN_t(WX7255_t),
    .SDIN(n7555),
    .SDIN_t(n7555_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7556),
    .Q_t(n7556_t),
    .QN(n5427),
    .QN_t(n5427_t)
  );


  sdffs1
  \DFF_1064/Q_reg 
  (
    .DIN(WX7253),
    .DIN_t(WX7253_t),
    .SDIN(n7554),
    .SDIN_t(n7554_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7555),
    .Q_t(n7555_t),
    .QN(n5432),
    .QN_t(n5432_t)
  );


  sdffs1
  \DFF_1063/Q_reg 
  (
    .DIN(WX7251),
    .DIN_t(WX7251_t),
    .SDIN(n7553),
    .SDIN_t(n7553_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7554),
    .Q_t(n7554_t),
    .QN(n5437),
    .QN_t(n5437_t)
  );


  sdffs1
  \DFF_1062/Q_reg 
  (
    .DIN(WX7249),
    .DIN_t(WX7249_t),
    .SDIN(n7552),
    .SDIN_t(n7552_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7553),
    .Q_t(n7553_t),
    .QN(n5442),
    .QN_t(n5442_t)
  );


  sdffs1
  \DFF_1061/Q_reg 
  (
    .DIN(WX7247),
    .DIN_t(WX7247_t),
    .SDIN(n7551),
    .SDIN_t(n7551_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7552),
    .Q_t(n7552_t),
    .QN(n5447),
    .QN_t(n5447_t)
  );


  sdffs1
  \DFF_1060/Q_reg 
  (
    .DIN(WX7245),
    .DIN_t(WX7245_t),
    .SDIN(n7550),
    .SDIN_t(n7550_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7551),
    .Q_t(n7551_t),
    .QN(n5452),
    .QN_t(n5452_t)
  );


  sdffs1
  \DFF_1059/Q_reg 
  (
    .DIN(WX7243),
    .DIN_t(WX7243_t),
    .SDIN(n7549),
    .SDIN_t(n7549_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7550),
    .Q_t(n7550_t),
    .QN(n5457),
    .QN_t(n5457_t)
  );


  sdffs1
  \DFF_1058/Q_reg 
  (
    .DIN(WX7241),
    .DIN_t(WX7241_t),
    .SDIN(n7548),
    .SDIN_t(n7548_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7549),
    .Q_t(n7549_t),
    .QN(n5462),
    .QN_t(n5462_t)
  );


  sdffs1
  \DFF_1057/Q_reg 
  (
    .DIN(WX7239),
    .DIN_t(WX7239_t),
    .SDIN(n7547),
    .SDIN_t(n7547_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7548),
    .Q_t(n7548_t),
    .QN(n5467),
    .QN_t(n5467_t)
  );


  sdffs1
  \DFF_1056/Q_reg 
  (
    .DIN(WX7237),
    .DIN_t(WX7237_t),
    .SDIN(n7546),
    .SDIN_t(n7546_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7547),
    .Q_t(n7547_t),
    .QN(n5472),
    .QN_t(n5472_t)
  );


  sdffs1
  \DFF_1055/Q_reg 
  (
    .DIN(WX7235),
    .DIN_t(WX7235_t),
    .SDIN(n7545),
    .SDIN_t(n7545_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7546),
    .Q_t(n7546_t),
    .QN(n5332),
    .QN_t(n5332_t)
  );


  sdffs1
  \DFF_1054/Q_reg 
  (
    .DIN(WX7233),
    .DIN_t(WX7233_t),
    .SDIN(n7544),
    .SDIN_t(n7544_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7545),
    .Q_t(n7545_t),
    .QN(n5336),
    .QN_t(n5336_t)
  );


  sdffs1
  \DFF_1053/Q_reg 
  (
    .DIN(WX7231),
    .DIN_t(WX7231_t),
    .SDIN(n7543),
    .SDIN_t(n7543_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7544),
    .Q_t(n7544_t),
    .QN(n5340),
    .QN_t(n5340_t)
  );


  sdffs1
  \DFF_1052/Q_reg 
  (
    .DIN(WX7229),
    .DIN_t(WX7229_t),
    .SDIN(n7542),
    .SDIN_t(n7542_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7543),
    .Q_t(n7543_t),
    .QN(n5344),
    .QN_t(n5344_t)
  );


  sdffs1
  \DFF_1051/Q_reg 
  (
    .DIN(WX7227),
    .DIN_t(WX7227_t),
    .SDIN(n7541),
    .SDIN_t(n7541_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7542),
    .Q_t(n7542_t),
    .QN(n5348),
    .QN_t(n5348_t)
  );


  sdffs1
  \DFF_1050/Q_reg 
  (
    .DIN(WX7225),
    .DIN_t(WX7225_t),
    .SDIN(n7540),
    .SDIN_t(n7540_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7541),
    .Q_t(n7541_t),
    .QN(n5352),
    .QN_t(n5352_t)
  );


  sdffs1
  \DFF_1049/Q_reg 
  (
    .DIN(WX7223),
    .DIN_t(WX7223_t),
    .SDIN(n7539),
    .SDIN_t(n7539_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7540),
    .Q_t(n7540_t),
    .QN(n5356),
    .QN_t(n5356_t)
  );


  sdffs1
  \DFF_1048/Q_reg 
  (
    .DIN(WX7221),
    .DIN_t(WX7221_t),
    .SDIN(n7538),
    .SDIN_t(n7538_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7539),
    .Q_t(n7539_t),
    .QN(n5360),
    .QN_t(n5360_t)
  );


  sdffs1
  \DFF_1047/Q_reg 
  (
    .DIN(WX7219),
    .DIN_t(WX7219_t),
    .SDIN(n7537),
    .SDIN_t(n7537_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7538),
    .Q_t(n7538_t),
    .QN(n5364),
    .QN_t(n5364_t)
  );


  sdffs1
  \DFF_1046/Q_reg 
  (
    .DIN(WX7217),
    .DIN_t(WX7217_t),
    .SDIN(n7536),
    .SDIN_t(n7536_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7537),
    .Q_t(n7537_t),
    .QN(n5368),
    .QN_t(n5368_t)
  );


  sdffs1
  \DFF_1045/Q_reg 
  (
    .DIN(WX7215),
    .DIN_t(WX7215_t),
    .SDIN(n7535),
    .SDIN_t(n7535_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7536),
    .Q_t(n7536_t),
    .QN(n5372),
    .QN_t(n5372_t)
  );


  sdffs1
  \DFF_1044/Q_reg 
  (
    .DIN(WX7213),
    .DIN_t(WX7213_t),
    .SDIN(n7534),
    .SDIN_t(n7534_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7535),
    .Q_t(n7535_t),
    .QN(n5376),
    .QN_t(n5376_t)
  );


  sdffs1
  \DFF_1043/Q_reg 
  (
    .DIN(WX7211),
    .DIN_t(WX7211_t),
    .SDIN(n7533),
    .SDIN_t(n7533_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7534),
    .Q_t(n7534_t),
    .QN(n5380),
    .QN_t(n5380_t)
  );


  sdffs1
  \DFF_1042/Q_reg 
  (
    .DIN(WX7209),
    .DIN_t(WX7209_t),
    .SDIN(n7532),
    .SDIN_t(n7532_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7533),
    .Q_t(n7533_t),
    .QN(n5384),
    .QN_t(n5384_t)
  );


  sdffs1
  \DFF_1041/Q_reg 
  (
    .DIN(WX7207),
    .DIN_t(WX7207_t),
    .SDIN(n7531),
    .SDIN_t(n7531_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7532),
    .Q_t(n7532_t),
    .QN(n5388),
    .QN_t(n5388_t)
  );


  sdffs1
  \DFF_1040/Q_reg 
  (
    .DIN(WX7205),
    .DIN_t(WX7205_t),
    .SDIN(n5396),
    .SDIN_t(n5396_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7531),
    .Q_t(n7531_t),
    .QN(n5392),
    .QN_t(n5392_t)
  );


  sdffs1
  \DFF_1039/Q_reg 
  (
    .DIN(WX7203),
    .DIN_t(WX7203_t),
    .SDIN(n5401),
    .SDIN_t(n5401_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5396),
    .Q_t(n5396_t)
  );


  sdffs1
  \DFF_1038/Q_reg 
  (
    .DIN(WX7201),
    .DIN_t(WX7201_t),
    .SDIN(n5406),
    .SDIN_t(n5406_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5401),
    .Q_t(n5401_t)
  );


  sdffs1
  \DFF_1037/Q_reg 
  (
    .DIN(WX7199),
    .DIN_t(WX7199_t),
    .SDIN(n5411),
    .SDIN_t(n5411_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5406),
    .Q_t(n5406_t)
  );


  sdffs1
  \DFF_1036/Q_reg 
  (
    .DIN(WX7197),
    .DIN_t(WX7197_t),
    .SDIN(n5416),
    .SDIN_t(n5416_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5411),
    .Q_t(n5411_t)
  );


  sdffs1
  \DFF_1035/Q_reg 
  (
    .DIN(WX7195),
    .DIN_t(WX7195_t),
    .SDIN(n5421),
    .SDIN_t(n5421_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5416),
    .Q_t(n5416_t)
  );


  sdffs1
  \DFF_1034/Q_reg 
  (
    .DIN(WX7193),
    .DIN_t(WX7193_t),
    .SDIN(n5426),
    .SDIN_t(n5426_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5421),
    .Q_t(n5421_t)
  );


  sdffs1
  \DFF_1033/Q_reg 
  (
    .DIN(WX7191),
    .DIN_t(WX7191_t),
    .SDIN(n5431),
    .SDIN_t(n5431_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5426),
    .Q_t(n5426_t)
  );


  sdffs1
  \DFF_1032/Q_reg 
  (
    .DIN(WX7189),
    .DIN_t(WX7189_t),
    .SDIN(n5436),
    .SDIN_t(n5436_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5431),
    .Q_t(n5431_t)
  );


  sdffs1
  \DFF_1031/Q_reg 
  (
    .DIN(WX7187),
    .DIN_t(WX7187_t),
    .SDIN(n5441),
    .SDIN_t(n5441_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5436),
    .Q_t(n5436_t)
  );


  sdffs1
  \DFF_1030/Q_reg 
  (
    .DIN(WX7185),
    .DIN_t(WX7185_t),
    .SDIN(n5446),
    .SDIN_t(n5446_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5441),
    .Q_t(n5441_t)
  );


  sdffs1
  \DFF_1029/Q_reg 
  (
    .DIN(WX7183),
    .DIN_t(WX7183_t),
    .SDIN(n5451),
    .SDIN_t(n5451_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5446),
    .Q_t(n5446_t)
  );


  sdffs1
  \DFF_1028/Q_reg 
  (
    .DIN(WX7181),
    .DIN_t(WX7181_t),
    .SDIN(n5456),
    .SDIN_t(n5456_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5451),
    .Q_t(n5451_t)
  );


  sdffs1
  \DFF_1027/Q_reg 
  (
    .DIN(WX7179),
    .DIN_t(WX7179_t),
    .SDIN(n5461),
    .SDIN_t(n5461_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5456),
    .Q_t(n5456_t)
  );


  sdffs1
  \DFF_1026/Q_reg 
  (
    .DIN(WX7177),
    .DIN_t(WX7177_t),
    .SDIN(n5466),
    .SDIN_t(n5466_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5461),
    .Q_t(n5461_t)
  );


  sdffs1
  \DFF_1025/Q_reg 
  (
    .DIN(WX7175),
    .DIN_t(WX7175_t),
    .SDIN(n5471),
    .SDIN_t(n5471_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5466),
    .Q_t(n5466_t)
  );


  sdffs1
  \DFF_1024/Q_reg 
  (
    .DIN(WX7173),
    .DIN_t(WX7173_t),
    .SDIN(n5331),
    .SDIN_t(n5331_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5471),
    .Q_t(n5471_t)
  );


  sdffs1
  \DFF_1023/Q_reg 
  (
    .DIN(WX7171),
    .DIN_t(WX7171_t),
    .SDIN(n5335),
    .SDIN_t(n5335_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5331),
    .Q_t(n5331_t)
  );


  sdffs1
  \DFF_1022/Q_reg 
  (
    .DIN(WX7169),
    .DIN_t(WX7169_t),
    .SDIN(n5339),
    .SDIN_t(n5339_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5335),
    .Q_t(n5335_t)
  );


  sdffs1
  \DFF_1021/Q_reg 
  (
    .DIN(WX7167),
    .DIN_t(WX7167_t),
    .SDIN(n5343),
    .SDIN_t(n5343_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5339),
    .Q_t(n5339_t)
  );


  sdffs1
  \DFF_1020/Q_reg 
  (
    .DIN(WX7165),
    .DIN_t(WX7165_t),
    .SDIN(n5347),
    .SDIN_t(n5347_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5343),
    .Q_t(n5343_t)
  );


  sdffs1
  \DFF_1019/Q_reg 
  (
    .DIN(WX7163),
    .DIN_t(WX7163_t),
    .SDIN(n5351),
    .SDIN_t(n5351_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5347),
    .Q_t(n5347_t)
  );


  sdffs1
  \DFF_1018/Q_reg 
  (
    .DIN(WX7161),
    .DIN_t(WX7161_t),
    .SDIN(n5355),
    .SDIN_t(n5355_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5351),
    .Q_t(n5351_t)
  );


  sdffs1
  \DFF_1017/Q_reg 
  (
    .DIN(WX7159),
    .DIN_t(WX7159_t),
    .SDIN(n5359),
    .SDIN_t(n5359_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5355),
    .Q_t(n5355_t)
  );


  sdffs1
  \DFF_1016/Q_reg 
  (
    .DIN(WX7157),
    .DIN_t(WX7157_t),
    .SDIN(n5363),
    .SDIN_t(n5363_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5359),
    .Q_t(n5359_t)
  );


  sdffs1
  \DFF_1015/Q_reg 
  (
    .DIN(WX7155),
    .DIN_t(WX7155_t),
    .SDIN(n5367),
    .SDIN_t(n5367_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5363),
    .Q_t(n5363_t)
  );


  sdffs1
  \DFF_1014/Q_reg 
  (
    .DIN(WX7153),
    .DIN_t(WX7153_t),
    .SDIN(n5371),
    .SDIN_t(n5371_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5367),
    .Q_t(n5367_t)
  );


  sdffs1
  \DFF_1013/Q_reg 
  (
    .DIN(WX7151),
    .DIN_t(WX7151_t),
    .SDIN(n5375),
    .SDIN_t(n5375_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5371),
    .Q_t(n5371_t)
  );


  sdffs1
  \DFF_1012/Q_reg 
  (
    .DIN(WX7149),
    .DIN_t(WX7149_t),
    .SDIN(n5379),
    .SDIN_t(n5379_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5375),
    .Q_t(n5375_t)
  );


  sdffs1
  \DFF_1011/Q_reg 
  (
    .DIN(WX7147),
    .DIN_t(WX7147_t),
    .SDIN(n5383),
    .SDIN_t(n5383_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5379),
    .Q_t(n5379_t)
  );


  sdffs1
  \DFF_1010/Q_reg 
  (
    .DIN(WX7145),
    .DIN_t(WX7145_t),
    .SDIN(n5387),
    .SDIN_t(n5387_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5383),
    .Q_t(n5383_t)
  );


  sdffs1
  \DFF_1009/Q_reg 
  (
    .DIN(WX7143),
    .DIN_t(WX7143_t),
    .SDIN(n5391),
    .SDIN_t(n5391_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5387),
    .Q_t(n5387_t)
  );


  sdffs1
  \DFF_1008/Q_reg 
  (
    .DIN(WX7141),
    .DIN_t(WX7141_t),
    .SDIN(n7530),
    .SDIN_t(n7530_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5391),
    .Q_t(n5391_t)
  );


  sdffs1
  \DFF_1007/Q_reg 
  (
    .DIN(WX7139),
    .DIN_t(WX7139_t),
    .SDIN(n7529),
    .SDIN_t(n7529_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7530),
    .Q_t(n7530_t),
    .QN(n5395),
    .QN_t(n5395_t)
  );


  sdffs1
  \DFF_1006/Q_reg 
  (
    .DIN(WX7137),
    .DIN_t(WX7137_t),
    .SDIN(n7528),
    .SDIN_t(n7528_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7529),
    .Q_t(n7529_t),
    .QN(n5400),
    .QN_t(n5400_t)
  );


  sdffs1
  \DFF_1005/Q_reg 
  (
    .DIN(WX7135),
    .DIN_t(WX7135_t),
    .SDIN(n7527),
    .SDIN_t(n7527_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7528),
    .Q_t(n7528_t),
    .QN(n5405),
    .QN_t(n5405_t)
  );


  sdffs1
  \DFF_1004/Q_reg 
  (
    .DIN(WX7133),
    .DIN_t(WX7133_t),
    .SDIN(n7526),
    .SDIN_t(n7526_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7527),
    .Q_t(n7527_t),
    .QN(n5410),
    .QN_t(n5410_t)
  );


  sdffs1
  \DFF_1003/Q_reg 
  (
    .DIN(WX7131),
    .DIN_t(WX7131_t),
    .SDIN(n7525),
    .SDIN_t(n7525_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7526),
    .Q_t(n7526_t),
    .QN(n5415),
    .QN_t(n5415_t)
  );


  sdffs1
  \DFF_1002/Q_reg 
  (
    .DIN(WX7129),
    .DIN_t(WX7129_t),
    .SDIN(n7524),
    .SDIN_t(n7524_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7525),
    .Q_t(n7525_t),
    .QN(n5420),
    .QN_t(n5420_t)
  );


  sdffs1
  \DFF_1001/Q_reg 
  (
    .DIN(WX7127),
    .DIN_t(WX7127_t),
    .SDIN(n7523),
    .SDIN_t(n7523_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7524),
    .Q_t(n7524_t),
    .QN(n5425),
    .QN_t(n5425_t)
  );


  sdffs1
  \DFF_1000/Q_reg 
  (
    .DIN(WX7125),
    .DIN_t(WX7125_t),
    .SDIN(n7522),
    .SDIN_t(n7522_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7523),
    .Q_t(n7523_t),
    .QN(n5430),
    .QN_t(n5430_t)
  );


  sdffs1
  \DFF_999/Q_reg 
  (
    .DIN(WX7123),
    .DIN_t(WX7123_t),
    .SDIN(n7521),
    .SDIN_t(n7521_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7522),
    .Q_t(n7522_t),
    .QN(n5435),
    .QN_t(n5435_t)
  );


  sdffs1
  \DFF_998/Q_reg 
  (
    .DIN(WX7121),
    .DIN_t(WX7121_t),
    .SDIN(n7520),
    .SDIN_t(n7520_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7521),
    .Q_t(n7521_t),
    .QN(n5440),
    .QN_t(n5440_t)
  );


  sdffs1
  \DFF_997/Q_reg 
  (
    .DIN(WX7119),
    .DIN_t(WX7119_t),
    .SDIN(n7519),
    .SDIN_t(n7519_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7520),
    .Q_t(n7520_t),
    .QN(n5445),
    .QN_t(n5445_t)
  );


  sdffs1
  \DFF_996/Q_reg 
  (
    .DIN(WX7117),
    .DIN_t(WX7117_t),
    .SDIN(n7518),
    .SDIN_t(n7518_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7519),
    .Q_t(n7519_t),
    .QN(n5450),
    .QN_t(n5450_t)
  );


  sdffs1
  \DFF_995/Q_reg 
  (
    .DIN(WX7115),
    .DIN_t(WX7115_t),
    .SDIN(n7517),
    .SDIN_t(n7517_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7518),
    .Q_t(n7518_t),
    .QN(n5455),
    .QN_t(n5455_t)
  );


  sdffs1
  \DFF_994/Q_reg 
  (
    .DIN(WX7113),
    .DIN_t(WX7113_t),
    .SDIN(n7516),
    .SDIN_t(n7516_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7517),
    .Q_t(n7517_t),
    .QN(n5460),
    .QN_t(n5460_t)
  );


  sdffs1
  \DFF_993/Q_reg 
  (
    .DIN(WX7111),
    .DIN_t(WX7111_t),
    .SDIN(n7515),
    .SDIN_t(n7515_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7516),
    .Q_t(n7516_t),
    .QN(n5465),
    .QN_t(n5465_t)
  );


  sdffs1
  \DFF_992/Q_reg 
  (
    .DIN(WX7109),
    .DIN_t(WX7109_t),
    .SDIN(n7514),
    .SDIN_t(n7514_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7515),
    .Q_t(n7515_t),
    .QN(n5470),
    .QN_t(n5470_t)
  );


  sdffs1
  \DFF_991/Q_reg 
  (
    .DIN(WX7011),
    .DIN_t(WX7011_t),
    .SDIN(n7513),
    .SDIN_t(n7513_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7514),
    .Q_t(n7514_t),
    .QN(n5300),
    .QN_t(n5300_t)
  );


  sdffs1
  \DFF_990/Q_reg 
  (
    .DIN(WX7009),
    .DIN_t(WX7009_t),
    .SDIN(n7512),
    .SDIN_t(n7512_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7513),
    .Q_t(n7513_t),
    .QN(n5301),
    .QN_t(n5301_t)
  );


  sdffs1
  \DFF_989/Q_reg 
  (
    .DIN(WX7007),
    .DIN_t(WX7007_t),
    .SDIN(n7511),
    .SDIN_t(n7511_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7512),
    .Q_t(n7512_t),
    .QN(n5302),
    .QN_t(n5302_t)
  );


  sdffs1
  \DFF_988/Q_reg 
  (
    .DIN(WX7005),
    .DIN_t(WX7005_t),
    .SDIN(n7510),
    .SDIN_t(n7510_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7511),
    .Q_t(n7511_t),
    .QN(n5303),
    .QN_t(n5303_t)
  );


  sdffs1
  \DFF_987/Q_reg 
  (
    .DIN(WX7003),
    .DIN_t(WX7003_t),
    .SDIN(n7509),
    .SDIN_t(n7509_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7510),
    .Q_t(n7510_t),
    .QN(n5304),
    .QN_t(n5304_t)
  );


  sdffs1
  \DFF_986/Q_reg 
  (
    .DIN(WX7001),
    .DIN_t(WX7001_t),
    .SDIN(n7508),
    .SDIN_t(n7508_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7509),
    .Q_t(n7509_t),
    .QN(n5305),
    .QN_t(n5305_t)
  );


  sdffs1
  \DFF_985/Q_reg 
  (
    .DIN(WX6999),
    .DIN_t(WX6999_t),
    .SDIN(n7507),
    .SDIN_t(n7507_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7508),
    .Q_t(n7508_t),
    .QN(n5306),
    .QN_t(n5306_t)
  );


  sdffs1
  \DFF_984/Q_reg 
  (
    .DIN(WX6997),
    .DIN_t(WX6997_t),
    .SDIN(n7506),
    .SDIN_t(n7506_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7507),
    .Q_t(n7507_t),
    .QN(n5307),
    .QN_t(n5307_t)
  );


  sdffs1
  \DFF_983/Q_reg 
  (
    .DIN(WX6995),
    .DIN_t(WX6995_t),
    .SDIN(n7505),
    .SDIN_t(n7505_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7506),
    .Q_t(n7506_t),
    .QN(n5308),
    .QN_t(n5308_t)
  );


  sdffs1
  \DFF_982/Q_reg 
  (
    .DIN(WX6993),
    .DIN_t(WX6993_t),
    .SDIN(n7504),
    .SDIN_t(n7504_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7505),
    .Q_t(n7505_t),
    .QN(n5309),
    .QN_t(n5309_t)
  );


  sdffs1
  \DFF_981/Q_reg 
  (
    .DIN(WX6991),
    .DIN_t(WX6991_t),
    .SDIN(n7503),
    .SDIN_t(n7503_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7504),
    .Q_t(n7504_t),
    .QN(n5310),
    .QN_t(n5310_t)
  );


  sdffs1
  \DFF_980/Q_reg 
  (
    .DIN(WX6989),
    .DIN_t(WX6989_t),
    .SDIN(n7502),
    .SDIN_t(n7502_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7503),
    .Q_t(n7503_t),
    .QN(n5311),
    .QN_t(n5311_t)
  );


  sdffs1
  \DFF_979/Q_reg 
  (
    .DIN(WX6987),
    .DIN_t(WX6987_t),
    .SDIN(n7501),
    .SDIN_t(n7501_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7502),
    .Q_t(n7502_t),
    .QN(n5312),
    .QN_t(n5312_t)
  );


  sdffs1
  \DFF_978/Q_reg 
  (
    .DIN(WX6985),
    .DIN_t(WX6985_t),
    .SDIN(n7500),
    .SDIN_t(n7500_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7501),
    .Q_t(n7501_t),
    .QN(n5313),
    .QN_t(n5313_t)
  );


  sdffs1
  \DFF_977/Q_reg 
  (
    .DIN(WX6983),
    .DIN_t(WX6983_t),
    .SDIN(n7499),
    .SDIN_t(n7499_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7500),
    .Q_t(n7500_t),
    .QN(n5314),
    .QN_t(n5314_t)
  );


  sdffs1
  \DFF_976/Q_reg 
  (
    .DIN(WX6981),
    .DIN_t(WX6981_t),
    .SDIN(n7498),
    .SDIN_t(n7498_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7499),
    .Q_t(n7499_t),
    .QN(n5315),
    .QN_t(n5315_t)
  );


  sdffs1
  \DFF_975/Q_reg 
  (
    .DIN(WX6979),
    .DIN_t(WX6979_t),
    .SDIN(n7497),
    .SDIN_t(n7497_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7498),
    .Q_t(n7498_t),
    .QN(n5316),
    .QN_t(n5316_t)
  );


  sdffs1
  \DFF_974/Q_reg 
  (
    .DIN(WX6977),
    .DIN_t(WX6977_t),
    .SDIN(n7496),
    .SDIN_t(n7496_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7497),
    .Q_t(n7497_t),
    .QN(n5317),
    .QN_t(n5317_t)
  );


  sdffs1
  \DFF_973/Q_reg 
  (
    .DIN(WX6975),
    .DIN_t(WX6975_t),
    .SDIN(n7495),
    .SDIN_t(n7495_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7496),
    .Q_t(n7496_t),
    .QN(n5318),
    .QN_t(n5318_t)
  );


  sdffs1
  \DFF_972/Q_reg 
  (
    .DIN(WX6973),
    .DIN_t(WX6973_t),
    .SDIN(n7494),
    .SDIN_t(n7494_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7495),
    .Q_t(n7495_t),
    .QN(n5319),
    .QN_t(n5319_t)
  );


  sdffs1
  \DFF_971/Q_reg 
  (
    .DIN(WX6971),
    .DIN_t(WX6971_t),
    .SDIN(n7493),
    .SDIN_t(n7493_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7494),
    .Q_t(n7494_t),
    .QN(n5320),
    .QN_t(n5320_t)
  );


  sdffs1
  \DFF_970/Q_reg 
  (
    .DIN(WX6969),
    .DIN_t(WX6969_t),
    .SDIN(n7492),
    .SDIN_t(n7492_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7493),
    .Q_t(n7493_t),
    .QN(n5321),
    .QN_t(n5321_t)
  );


  sdffs1
  \DFF_969/Q_reg 
  (
    .DIN(WX6967),
    .DIN_t(WX6967_t),
    .SDIN(n7491),
    .SDIN_t(n7491_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7492),
    .Q_t(n7492_t),
    .QN(n5322),
    .QN_t(n5322_t)
  );


  sdffs1
  \DFF_968/Q_reg 
  (
    .DIN(WX6965),
    .DIN_t(WX6965_t),
    .SDIN(n7490),
    .SDIN_t(n7490_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7491),
    .Q_t(n7491_t),
    .QN(n5323),
    .QN_t(n5323_t)
  );


  sdffs1
  \DFF_967/Q_reg 
  (
    .DIN(WX6963),
    .DIN_t(WX6963_t),
    .SDIN(n7489),
    .SDIN_t(n7489_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7490),
    .Q_t(n7490_t),
    .QN(n5324),
    .QN_t(n5324_t)
  );


  sdffs1
  \DFF_966/Q_reg 
  (
    .DIN(WX6961),
    .DIN_t(WX6961_t),
    .SDIN(n7488),
    .SDIN_t(n7488_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7489),
    .Q_t(n7489_t),
    .QN(n5325),
    .QN_t(n5325_t)
  );


  sdffs1
  \DFF_965/Q_reg 
  (
    .DIN(WX6959),
    .DIN_t(WX6959_t),
    .SDIN(n7487),
    .SDIN_t(n7487_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7488),
    .Q_t(n7488_t),
    .QN(n5326),
    .QN_t(n5326_t)
  );


  sdffs1
  \DFF_964/Q_reg 
  (
    .DIN(WX6957),
    .DIN_t(WX6957_t),
    .SDIN(n7486),
    .SDIN_t(n7486_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7487),
    .Q_t(n7487_t),
    .QN(n5327),
    .QN_t(n5327_t)
  );


  sdffs1
  \DFF_963/Q_reg 
  (
    .DIN(WX6955),
    .DIN_t(WX6955_t),
    .SDIN(n7485),
    .SDIN_t(n7485_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7486),
    .Q_t(n7486_t),
    .QN(n5328),
    .QN_t(n5328_t)
  );


  sdffs1
  \DFF_962/Q_reg 
  (
    .DIN(WX6953),
    .DIN_t(WX6953_t),
    .SDIN(n7484),
    .SDIN_t(n7484_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7485),
    .Q_t(n7485_t),
    .QN(n5329),
    .QN_t(n5329_t)
  );


  sdffs1
  \DFF_961/Q_reg 
  (
    .DIN(WX6951),
    .DIN_t(WX6951_t),
    .SDIN(n7483),
    .SDIN_t(n7483_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7484),
    .Q_t(n7484_t),
    .QN(n5330),
    .QN_t(n5330_t)
  );


  sdffs1
  \DFF_960/Q_reg 
  (
    .DIN(WX6949),
    .DIN_t(WX6949_t),
    .SDIN(CRC_OUT_5_31),
    .SDIN_t(CRC_OUT_5_31_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7483),
    .Q_t(n7483_t),
    .QN(n5299),
    .QN_t(n5299_t)
  );


  sdffs1
  \DFF_959/Q_reg 
  (
    .DIN(WX6498),
    .DIN_t(WX6498_t),
    .SDIN(CRC_OUT_5_30),
    .SDIN_t(CRC_OUT_5_30_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_31),
    .Q_t(CRC_OUT_5_31_t),
    .QN(n5474),
    .QN_t(n5474_t)
  );


  sdffs1
  \DFF_958/Q_reg 
  (
    .DIN(WX6496),
    .DIN_t(WX6496_t),
    .SDIN(CRC_OUT_5_29),
    .SDIN_t(CRC_OUT_5_29_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_30),
    .Q_t(CRC_OUT_5_30_t),
    .QN(n5469),
    .QN_t(n5469_t)
  );


  sdffs1
  \DFF_957/Q_reg 
  (
    .DIN(WX6494),
    .DIN_t(WX6494_t),
    .SDIN(CRC_OUT_5_28),
    .SDIN_t(CRC_OUT_5_28_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_29),
    .Q_t(CRC_OUT_5_29_t),
    .QN(n5464),
    .QN_t(n5464_t)
  );


  sdffs1
  \DFF_956/Q_reg 
  (
    .DIN(WX6492),
    .DIN_t(WX6492_t),
    .SDIN(CRC_OUT_5_27),
    .SDIN_t(CRC_OUT_5_27_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_28),
    .Q_t(CRC_OUT_5_28_t),
    .QN(n5459),
    .QN_t(n5459_t)
  );


  sdffs1
  \DFF_955/Q_reg 
  (
    .DIN(WX6490),
    .DIN_t(WX6490_t),
    .SDIN(CRC_OUT_5_26),
    .SDIN_t(CRC_OUT_5_26_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_27),
    .Q_t(CRC_OUT_5_27_t),
    .QN(n5454),
    .QN_t(n5454_t)
  );


  sdffs1
  \DFF_954/Q_reg 
  (
    .DIN(WX6488),
    .DIN_t(WX6488_t),
    .SDIN(CRC_OUT_5_25),
    .SDIN_t(CRC_OUT_5_25_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_26),
    .Q_t(CRC_OUT_5_26_t),
    .QN(n5449),
    .QN_t(n5449_t)
  );


  sdffs1
  \DFF_953/Q_reg 
  (
    .DIN(WX6486),
    .DIN_t(WX6486_t),
    .SDIN(CRC_OUT_5_24),
    .SDIN_t(CRC_OUT_5_24_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_25),
    .Q_t(CRC_OUT_5_25_t),
    .QN(n5444),
    .QN_t(n5444_t)
  );


  sdffs1
  \DFF_952/Q_reg 
  (
    .DIN(WX6484),
    .DIN_t(WX6484_t),
    .SDIN(CRC_OUT_5_23),
    .SDIN_t(CRC_OUT_5_23_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_24),
    .Q_t(CRC_OUT_5_24_t),
    .QN(n5439),
    .QN_t(n5439_t)
  );


  sdffs1
  \DFF_951/Q_reg 
  (
    .DIN(WX6482),
    .DIN_t(WX6482_t),
    .SDIN(CRC_OUT_5_22),
    .SDIN_t(CRC_OUT_5_22_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_23),
    .Q_t(CRC_OUT_5_23_t),
    .QN(n5434),
    .QN_t(n5434_t)
  );


  sdffs1
  \DFF_950/Q_reg 
  (
    .DIN(WX6480),
    .DIN_t(WX6480_t),
    .SDIN(CRC_OUT_5_21),
    .SDIN_t(CRC_OUT_5_21_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_22),
    .Q_t(CRC_OUT_5_22_t),
    .QN(n5429),
    .QN_t(n5429_t)
  );


  sdffs1
  \DFF_949/Q_reg 
  (
    .DIN(WX6478),
    .DIN_t(WX6478_t),
    .SDIN(CRC_OUT_5_20),
    .SDIN_t(CRC_OUT_5_20_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_21),
    .Q_t(CRC_OUT_5_21_t),
    .QN(n5424),
    .QN_t(n5424_t)
  );


  sdffs1
  \DFF_948/Q_reg 
  (
    .DIN(WX6476),
    .DIN_t(WX6476_t),
    .SDIN(CRC_OUT_5_19),
    .SDIN_t(CRC_OUT_5_19_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_20),
    .Q_t(CRC_OUT_5_20_t),
    .QN(n5419),
    .QN_t(n5419_t)
  );


  sdffs1
  \DFF_947/Q_reg 
  (
    .DIN(WX6474),
    .DIN_t(WX6474_t),
    .SDIN(CRC_OUT_5_18),
    .SDIN_t(CRC_OUT_5_18_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_19),
    .Q_t(CRC_OUT_5_19_t),
    .QN(n5414),
    .QN_t(n5414_t)
  );


  sdffs1
  \DFF_946/Q_reg 
  (
    .DIN(WX6472),
    .DIN_t(WX6472_t),
    .SDIN(CRC_OUT_5_17),
    .SDIN_t(CRC_OUT_5_17_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_18),
    .Q_t(CRC_OUT_5_18_t),
    .QN(n5409),
    .QN_t(n5409_t)
  );


  sdffs1
  \DFF_945/Q_reg 
  (
    .DIN(WX6470),
    .DIN_t(WX6470_t),
    .SDIN(CRC_OUT_5_16),
    .SDIN_t(CRC_OUT_5_16_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_17),
    .Q_t(CRC_OUT_5_17_t),
    .QN(n5404),
    .QN_t(n5404_t)
  );


  sdffs1
  \DFF_944/Q_reg 
  (
    .DIN(WX6468),
    .DIN_t(WX6468_t),
    .SDIN(CRC_OUT_5_15),
    .SDIN_t(CRC_OUT_5_15_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_16),
    .Q_t(CRC_OUT_5_16_t),
    .QN(n5399),
    .QN_t(n5399_t)
  );


  sdffs1
  \DFF_943/Q_reg 
  (
    .DIN(WX6466),
    .DIN_t(WX6466_t),
    .SDIN(CRC_OUT_5_14),
    .SDIN_t(CRC_OUT_5_14_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_15),
    .Q_t(CRC_OUT_5_15_t),
    .QN(n5394),
    .QN_t(n5394_t)
  );


  sdffs1
  \DFF_942/Q_reg 
  (
    .DIN(WX6464),
    .DIN_t(WX6464_t),
    .SDIN(CRC_OUT_5_13),
    .SDIN_t(CRC_OUT_5_13_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_14),
    .Q_t(CRC_OUT_5_14_t),
    .QN(n5390),
    .QN_t(n5390_t)
  );


  sdffs1
  \DFF_941/Q_reg 
  (
    .DIN(WX6462),
    .DIN_t(WX6462_t),
    .SDIN(CRC_OUT_5_12),
    .SDIN_t(CRC_OUT_5_12_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_13),
    .Q_t(CRC_OUT_5_13_t),
    .QN(n5386),
    .QN_t(n5386_t)
  );


  sdffs1
  \DFF_940/Q_reg 
  (
    .DIN(WX6460),
    .DIN_t(WX6460_t),
    .SDIN(CRC_OUT_5_11),
    .SDIN_t(CRC_OUT_5_11_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_12),
    .Q_t(CRC_OUT_5_12_t),
    .QN(n5382),
    .QN_t(n5382_t)
  );


  sdffs1
  \DFF_939/Q_reg 
  (
    .DIN(WX6458),
    .DIN_t(WX6458_t),
    .SDIN(CRC_OUT_5_10),
    .SDIN_t(CRC_OUT_5_10_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_11),
    .Q_t(CRC_OUT_5_11_t),
    .QN(n5378),
    .QN_t(n5378_t)
  );


  sdffs1
  \DFF_938/Q_reg 
  (
    .DIN(WX6456),
    .DIN_t(WX6456_t),
    .SDIN(CRC_OUT_5_9),
    .SDIN_t(CRC_OUT_5_9_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_10),
    .Q_t(CRC_OUT_5_10_t),
    .QN(n5374),
    .QN_t(n5374_t)
  );


  sdffs1
  \DFF_937/Q_reg 
  (
    .DIN(WX6454),
    .DIN_t(WX6454_t),
    .SDIN(CRC_OUT_5_8),
    .SDIN_t(CRC_OUT_5_8_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_9),
    .Q_t(CRC_OUT_5_9_t),
    .QN(n5370),
    .QN_t(n5370_t)
  );


  sdffs1
  \DFF_936/Q_reg 
  (
    .DIN(WX6452),
    .DIN_t(WX6452_t),
    .SDIN(CRC_OUT_5_7),
    .SDIN_t(CRC_OUT_5_7_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_8),
    .Q_t(CRC_OUT_5_8_t),
    .QN(n5366),
    .QN_t(n5366_t)
  );


  sdffs1
  \DFF_935/Q_reg 
  (
    .DIN(WX6450),
    .DIN_t(WX6450_t),
    .SDIN(CRC_OUT_5_6),
    .SDIN_t(CRC_OUT_5_6_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_7),
    .Q_t(CRC_OUT_5_7_t),
    .QN(n5362),
    .QN_t(n5362_t)
  );


  sdffs1
  \DFF_934/Q_reg 
  (
    .DIN(WX6448),
    .DIN_t(WX6448_t),
    .SDIN(CRC_OUT_5_5),
    .SDIN_t(CRC_OUT_5_5_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_6),
    .Q_t(CRC_OUT_5_6_t),
    .QN(n5358),
    .QN_t(n5358_t)
  );


  sdffs1
  \DFF_933/Q_reg 
  (
    .DIN(WX6446),
    .DIN_t(WX6446_t),
    .SDIN(CRC_OUT_5_4),
    .SDIN_t(CRC_OUT_5_4_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_5),
    .Q_t(CRC_OUT_5_5_t),
    .QN(n5354),
    .QN_t(n5354_t)
  );


  sdffs1
  \DFF_932/Q_reg 
  (
    .DIN(WX6444),
    .DIN_t(WX6444_t),
    .SDIN(CRC_OUT_5_3),
    .SDIN_t(CRC_OUT_5_3_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_4),
    .Q_t(CRC_OUT_5_4_t),
    .QN(n5350),
    .QN_t(n5350_t)
  );


  sdffs1
  \DFF_931/Q_reg 
  (
    .DIN(WX6442),
    .DIN_t(WX6442_t),
    .SDIN(CRC_OUT_5_2),
    .SDIN_t(CRC_OUT_5_2_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_3),
    .Q_t(CRC_OUT_5_3_t),
    .QN(n5346),
    .QN_t(n5346_t)
  );


  sdffs1
  \DFF_930/Q_reg 
  (
    .DIN(WX6440),
    .DIN_t(WX6440_t),
    .SDIN(CRC_OUT_5_1),
    .SDIN_t(CRC_OUT_5_1_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_2),
    .Q_t(CRC_OUT_5_2_t),
    .QN(n5342),
    .QN_t(n5342_t)
  );


  sdffs1
  \DFF_929/Q_reg 
  (
    .DIN(WX6438),
    .DIN_t(WX6438_t),
    .SDIN(CRC_OUT_5_0),
    .SDIN_t(CRC_OUT_5_0_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_1),
    .Q_t(CRC_OUT_5_1_t),
    .QN(n5338),
    .QN_t(n5338_t)
  );


  sdffs1
  \DFF_928/Q_reg 
  (
    .DIN(WX6436),
    .DIN_t(WX6436_t),
    .SDIN(n7482),
    .SDIN_t(n7482_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_5_0),
    .Q_t(CRC_OUT_5_0_t),
    .QN(n5334),
    .QN_t(n5334_t)
  );


  sdffs1
  \DFF_927/Q_reg 
  (
    .DIN(WX6070),
    .DIN_t(WX6070_t),
    .SDIN(n7481),
    .SDIN_t(n7481_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7482),
    .Q_t(n7482_t),
    .QN(n3253),
    .QN_t(n3253_t)
  );


  sdffs1
  \DFF_926/Q_reg 
  (
    .DIN(WX6068),
    .DIN_t(WX6068_t),
    .SDIN(n7480),
    .SDIN_t(n7480_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7481),
    .Q_t(n7481_t),
    .QN(n3254),
    .QN_t(n3254_t)
  );


  sdffs1
  \DFF_925/Q_reg 
  (
    .DIN(WX6066),
    .DIN_t(WX6066_t),
    .SDIN(n7479),
    .SDIN_t(n7479_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7480),
    .Q_t(n7480_t),
    .QN(n3255),
    .QN_t(n3255_t)
  );


  sdffs1
  \DFF_924/Q_reg 
  (
    .DIN(WX6064),
    .DIN_t(WX6064_t),
    .SDIN(n7478),
    .SDIN_t(n7478_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7479),
    .Q_t(n7479_t),
    .QN(n3256),
    .QN_t(n3256_t)
  );


  sdffs1
  \DFF_923/Q_reg 
  (
    .DIN(WX6062),
    .DIN_t(WX6062_t),
    .SDIN(n7477),
    .SDIN_t(n7477_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7478),
    .Q_t(n7478_t),
    .QN(n3257),
    .QN_t(n3257_t)
  );


  sdffs1
  \DFF_922/Q_reg 
  (
    .DIN(WX6060),
    .DIN_t(WX6060_t),
    .SDIN(n7476),
    .SDIN_t(n7476_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7477),
    .Q_t(n7477_t),
    .QN(n3258),
    .QN_t(n3258_t)
  );


  sdffs1
  \DFF_921/Q_reg 
  (
    .DIN(WX6058),
    .DIN_t(WX6058_t),
    .SDIN(n7475),
    .SDIN_t(n7475_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7476),
    .Q_t(n7476_t),
    .QN(n3259),
    .QN_t(n3259_t)
  );


  sdffs1
  \DFF_920/Q_reg 
  (
    .DIN(WX6056),
    .DIN_t(WX6056_t),
    .SDIN(n7474),
    .SDIN_t(n7474_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7475),
    .Q_t(n7475_t),
    .QN(n3260),
    .QN_t(n3260_t)
  );


  sdffs1
  \DFF_919/Q_reg 
  (
    .DIN(WX6054),
    .DIN_t(WX6054_t),
    .SDIN(n7473),
    .SDIN_t(n7473_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7474),
    .Q_t(n7474_t),
    .QN(n3261),
    .QN_t(n3261_t)
  );


  sdffs1
  \DFF_918/Q_reg 
  (
    .DIN(WX6052),
    .DIN_t(WX6052_t),
    .SDIN(n7472),
    .SDIN_t(n7472_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7473),
    .Q_t(n7473_t),
    .QN(n3262),
    .QN_t(n3262_t)
  );


  sdffs1
  \DFF_917/Q_reg 
  (
    .DIN(WX6050),
    .DIN_t(WX6050_t),
    .SDIN(n7471),
    .SDIN_t(n7471_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7472),
    .Q_t(n7472_t),
    .QN(n3263),
    .QN_t(n3263_t)
  );


  sdffs1
  \DFF_916/Q_reg 
  (
    .DIN(WX6048),
    .DIN_t(WX6048_t),
    .SDIN(n7470),
    .SDIN_t(n7470_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7471),
    .Q_t(n7471_t),
    .QN(n3264),
    .QN_t(n3264_t)
  );


  sdffs1
  \DFF_915/Q_reg 
  (
    .DIN(WX6046),
    .DIN_t(WX6046_t),
    .SDIN(n7469),
    .SDIN_t(n7469_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7470),
    .Q_t(n7470_t),
    .QN(n3265),
    .QN_t(n3265_t)
  );


  sdffs1
  \DFF_914/Q_reg 
  (
    .DIN(WX6044),
    .DIN_t(WX6044_t),
    .SDIN(n7468),
    .SDIN_t(n7468_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7469),
    .Q_t(n7469_t),
    .QN(n3266),
    .QN_t(n3266_t)
  );


  sdffs1
  \DFF_913/Q_reg 
  (
    .DIN(WX6042),
    .DIN_t(WX6042_t),
    .SDIN(n7467),
    .SDIN_t(n7467_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7468),
    .Q_t(n7468_t),
    .QN(n3267),
    .QN_t(n3267_t)
  );


  sdffs1
  \DFF_912/Q_reg 
  (
    .DIN(WX6040),
    .DIN_t(WX6040_t),
    .SDIN(n7466),
    .SDIN_t(n7466_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7467),
    .Q_t(n7467_t),
    .QN(n3268),
    .QN_t(n3268_t)
  );


  sdffs1
  \DFF_911/Q_reg 
  (
    .DIN(WX6038),
    .DIN_t(WX6038_t),
    .SDIN(n7465),
    .SDIN_t(n7465_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7466),
    .Q_t(n7466_t),
    .QN(n5574),
    .QN_t(n5574_t)
  );


  sdffs1
  \DFF_910/Q_reg 
  (
    .DIN(WX6036),
    .DIN_t(WX6036_t),
    .SDIN(n7464),
    .SDIN_t(n7464_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7465),
    .Q_t(n7465_t),
    .QN(n5579),
    .QN_t(n5579_t)
  );


  sdffs1
  \DFF_909/Q_reg 
  (
    .DIN(WX6034),
    .DIN_t(WX6034_t),
    .SDIN(n7463),
    .SDIN_t(n7463_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7464),
    .Q_t(n7464_t),
    .QN(n5584),
    .QN_t(n5584_t)
  );


  sdffs1
  \DFF_908/Q_reg 
  (
    .DIN(WX6032),
    .DIN_t(WX6032_t),
    .SDIN(n7462),
    .SDIN_t(n7462_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7463),
    .Q_t(n7463_t),
    .QN(n5589),
    .QN_t(n5589_t)
  );


  sdffs1
  \DFF_907/Q_reg 
  (
    .DIN(WX6030),
    .DIN_t(WX6030_t),
    .SDIN(n7461),
    .SDIN_t(n7461_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7462),
    .Q_t(n7462_t),
    .QN(n5594),
    .QN_t(n5594_t)
  );


  sdffs1
  \DFF_906/Q_reg 
  (
    .DIN(WX6028),
    .DIN_t(WX6028_t),
    .SDIN(n7460),
    .SDIN_t(n7460_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7461),
    .Q_t(n7461_t),
    .QN(n5599),
    .QN_t(n5599_t)
  );


  sdffs1
  \DFF_905/Q_reg 
  (
    .DIN(WX6026),
    .DIN_t(WX6026_t),
    .SDIN(n7459),
    .SDIN_t(n7459_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7460),
    .Q_t(n7460_t),
    .QN(n5604),
    .QN_t(n5604_t)
  );


  sdffs1
  \DFF_904/Q_reg 
  (
    .DIN(WX6024),
    .DIN_t(WX6024_t),
    .SDIN(n7458),
    .SDIN_t(n7458_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7459),
    .Q_t(n7459_t),
    .QN(n5609),
    .QN_t(n5609_t)
  );


  sdffs1
  \DFF_903/Q_reg 
  (
    .DIN(WX6022),
    .DIN_t(WX6022_t),
    .SDIN(n7457),
    .SDIN_t(n7457_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7458),
    .Q_t(n7458_t),
    .QN(n5614),
    .QN_t(n5614_t)
  );


  sdffs1
  \DFF_902/Q_reg 
  (
    .DIN(WX6020),
    .DIN_t(WX6020_t),
    .SDIN(n7456),
    .SDIN_t(n7456_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7457),
    .Q_t(n7457_t),
    .QN(n5619),
    .QN_t(n5619_t)
  );


  sdffs1
  \DFF_901/Q_reg 
  (
    .DIN(WX6018),
    .DIN_t(WX6018_t),
    .SDIN(n7455),
    .SDIN_t(n7455_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7456),
    .Q_t(n7456_t),
    .QN(n5624),
    .QN_t(n5624_t)
  );


  sdffs1
  \DFF_900/Q_reg 
  (
    .DIN(WX6016),
    .DIN_t(WX6016_t),
    .SDIN(n7454),
    .SDIN_t(n7454_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7455),
    .Q_t(n7455_t),
    .QN(n5629),
    .QN_t(n5629_t)
  );


  sdffs1
  \DFF_899/Q_reg 
  (
    .DIN(WX6014),
    .DIN_t(WX6014_t),
    .SDIN(n7453),
    .SDIN_t(n7453_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7454),
    .Q_t(n7454_t),
    .QN(n5634),
    .QN_t(n5634_t)
  );


  sdffs1
  \DFF_898/Q_reg 
  (
    .DIN(WX6012),
    .DIN_t(WX6012_t),
    .SDIN(n7452),
    .SDIN_t(n7452_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7453),
    .Q_t(n7453_t),
    .QN(n5639),
    .QN_t(n5639_t)
  );


  sdffs1
  \DFF_897/Q_reg 
  (
    .DIN(WX6010),
    .DIN_t(WX6010_t),
    .SDIN(n7451),
    .SDIN_t(n7451_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7452),
    .Q_t(n7452_t),
    .QN(n5644),
    .QN_t(n5644_t)
  );


  sdffs1
  \DFF_896/Q_reg 
  (
    .DIN(WX6008),
    .DIN_t(WX6008_t),
    .SDIN(n7450),
    .SDIN_t(n7450_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7451),
    .Q_t(n7451_t),
    .QN(n5649),
    .QN_t(n5649_t)
  );


  sdffs1
  \DFF_895/Q_reg 
  (
    .DIN(WX6006),
    .DIN_t(WX6006_t),
    .SDIN(n7449),
    .SDIN_t(n7449_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7450),
    .Q_t(n7450_t),
    .QN(n5509),
    .QN_t(n5509_t)
  );


  sdffs1
  \DFF_894/Q_reg 
  (
    .DIN(WX6004),
    .DIN_t(WX6004_t),
    .SDIN(n7448),
    .SDIN_t(n7448_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7449),
    .Q_t(n7449_t),
    .QN(n5513),
    .QN_t(n5513_t)
  );


  sdffs1
  \DFF_893/Q_reg 
  (
    .DIN(WX6002),
    .DIN_t(WX6002_t),
    .SDIN(n7447),
    .SDIN_t(n7447_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7448),
    .Q_t(n7448_t),
    .QN(n5517),
    .QN_t(n5517_t)
  );


  sdffs1
  \DFF_892/Q_reg 
  (
    .DIN(WX6000),
    .DIN_t(WX6000_t),
    .SDIN(n7446),
    .SDIN_t(n7446_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7447),
    .Q_t(n7447_t),
    .QN(n5521),
    .QN_t(n5521_t)
  );


  sdffs1
  \DFF_891/Q_reg 
  (
    .DIN(WX5998),
    .DIN_t(WX5998_t),
    .SDIN(n7445),
    .SDIN_t(n7445_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7446),
    .Q_t(n7446_t),
    .QN(n5525),
    .QN_t(n5525_t)
  );


  sdffs1
  \DFF_890/Q_reg 
  (
    .DIN(WX5996),
    .DIN_t(WX5996_t),
    .SDIN(n7444),
    .SDIN_t(n7444_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7445),
    .Q_t(n7445_t),
    .QN(n5529),
    .QN_t(n5529_t)
  );


  sdffs1
  \DFF_889/Q_reg 
  (
    .DIN(WX5994),
    .DIN_t(WX5994_t),
    .SDIN(n7443),
    .SDIN_t(n7443_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7444),
    .Q_t(n7444_t),
    .QN(n5533),
    .QN_t(n5533_t)
  );


  sdffs1
  \DFF_888/Q_reg 
  (
    .DIN(WX5992),
    .DIN_t(WX5992_t),
    .SDIN(n7442),
    .SDIN_t(n7442_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7443),
    .Q_t(n7443_t),
    .QN(n5537),
    .QN_t(n5537_t)
  );


  sdffs1
  \DFF_887/Q_reg 
  (
    .DIN(WX5990),
    .DIN_t(WX5990_t),
    .SDIN(n7441),
    .SDIN_t(n7441_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7442),
    .Q_t(n7442_t),
    .QN(n5541),
    .QN_t(n5541_t)
  );


  sdffs1
  \DFF_886/Q_reg 
  (
    .DIN(WX5988),
    .DIN_t(WX5988_t),
    .SDIN(n7440),
    .SDIN_t(n7440_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7441),
    .Q_t(n7441_t),
    .QN(n5545),
    .QN_t(n5545_t)
  );


  sdffs1
  \DFF_885/Q_reg 
  (
    .DIN(WX5986),
    .DIN_t(WX5986_t),
    .SDIN(n7439),
    .SDIN_t(n7439_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7440),
    .Q_t(n7440_t),
    .QN(n5549),
    .QN_t(n5549_t)
  );


  sdffs1
  \DFF_884/Q_reg 
  (
    .DIN(WX5984),
    .DIN_t(WX5984_t),
    .SDIN(n7438),
    .SDIN_t(n7438_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7439),
    .Q_t(n7439_t),
    .QN(n5553),
    .QN_t(n5553_t)
  );


  sdffs1
  \DFF_883/Q_reg 
  (
    .DIN(WX5982),
    .DIN_t(WX5982_t),
    .SDIN(n7437),
    .SDIN_t(n7437_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7438),
    .Q_t(n7438_t),
    .QN(n5557),
    .QN_t(n5557_t)
  );


  sdffs1
  \DFF_882/Q_reg 
  (
    .DIN(WX5980),
    .DIN_t(WX5980_t),
    .SDIN(n7436),
    .SDIN_t(n7436_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7437),
    .Q_t(n7437_t),
    .QN(n5561),
    .QN_t(n5561_t)
  );


  sdffs1
  \DFF_881/Q_reg 
  (
    .DIN(WX5978),
    .DIN_t(WX5978_t),
    .SDIN(n7435),
    .SDIN_t(n7435_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7436),
    .Q_t(n7436_t),
    .QN(n5565),
    .QN_t(n5565_t)
  );


  sdffs1
  \DFF_880/Q_reg 
  (
    .DIN(WX5976),
    .DIN_t(WX5976_t),
    .SDIN(n7434),
    .SDIN_t(n7434_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7435),
    .Q_t(n7435_t),
    .QN(n5569),
    .QN_t(n5569_t)
  );


  sdffs1
  \DFF_879/Q_reg 
  (
    .DIN(WX5974),
    .DIN_t(WX5974_t),
    .SDIN(n7433),
    .SDIN_t(n7433_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7434),
    .Q_t(n7434_t),
    .QN(n5573),
    .QN_t(n5573_t)
  );


  sdffs1
  \DFF_878/Q_reg 
  (
    .DIN(WX5972),
    .DIN_t(WX5972_t),
    .SDIN(n7432),
    .SDIN_t(n7432_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7433),
    .Q_t(n7433_t),
    .QN(n5578),
    .QN_t(n5578_t)
  );


  sdffs1
  \DFF_877/Q_reg 
  (
    .DIN(WX5970),
    .DIN_t(WX5970_t),
    .SDIN(n7431),
    .SDIN_t(n7431_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7432),
    .Q_t(n7432_t),
    .QN(n5583),
    .QN_t(n5583_t)
  );


  sdffs1
  \DFF_876/Q_reg 
  (
    .DIN(WX5968),
    .DIN_t(WX5968_t),
    .SDIN(n7430),
    .SDIN_t(n7430_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7431),
    .Q_t(n7431_t),
    .QN(n5588),
    .QN_t(n5588_t)
  );


  sdffs1
  \DFF_875/Q_reg 
  (
    .DIN(WX5966),
    .DIN_t(WX5966_t),
    .SDIN(n7429),
    .SDIN_t(n7429_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7430),
    .Q_t(n7430_t),
    .QN(n5593),
    .QN_t(n5593_t)
  );


  sdffs1
  \DFF_874/Q_reg 
  (
    .DIN(WX5964),
    .DIN_t(WX5964_t),
    .SDIN(n7428),
    .SDIN_t(n7428_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7429),
    .Q_t(n7429_t),
    .QN(n5598),
    .QN_t(n5598_t)
  );


  sdffs1
  \DFF_873/Q_reg 
  (
    .DIN(WX5962),
    .DIN_t(WX5962_t),
    .SDIN(n7427),
    .SDIN_t(n7427_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7428),
    .Q_t(n7428_t),
    .QN(n5603),
    .QN_t(n5603_t)
  );


  sdffs1
  \DFF_872/Q_reg 
  (
    .DIN(WX5960),
    .DIN_t(WX5960_t),
    .SDIN(n7426),
    .SDIN_t(n7426_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7427),
    .Q_t(n7427_t),
    .QN(n5608),
    .QN_t(n5608_t)
  );


  sdffs1
  \DFF_871/Q_reg 
  (
    .DIN(WX5958),
    .DIN_t(WX5958_t),
    .SDIN(n7425),
    .SDIN_t(n7425_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7426),
    .Q_t(n7426_t),
    .QN(n5613),
    .QN_t(n5613_t)
  );


  sdffs1
  \DFF_870/Q_reg 
  (
    .DIN(WX5956),
    .DIN_t(WX5956_t),
    .SDIN(n7424),
    .SDIN_t(n7424_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7425),
    .Q_t(n7425_t),
    .QN(n5618),
    .QN_t(n5618_t)
  );


  sdffs1
  \DFF_869/Q_reg 
  (
    .DIN(WX5954),
    .DIN_t(WX5954_t),
    .SDIN(n7423),
    .SDIN_t(n7423_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7424),
    .Q_t(n7424_t),
    .QN(n5623),
    .QN_t(n5623_t)
  );


  sdffs1
  \DFF_868/Q_reg 
  (
    .DIN(WX5952),
    .DIN_t(WX5952_t),
    .SDIN(n7422),
    .SDIN_t(n7422_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7423),
    .Q_t(n7423_t),
    .QN(n5628),
    .QN_t(n5628_t)
  );


  sdffs1
  \DFF_867/Q_reg 
  (
    .DIN(WX5950),
    .DIN_t(WX5950_t),
    .SDIN(n7421),
    .SDIN_t(n7421_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7422),
    .Q_t(n7422_t),
    .QN(n5633),
    .QN_t(n5633_t)
  );


  sdffs1
  \DFF_866/Q_reg 
  (
    .DIN(WX5948),
    .DIN_t(WX5948_t),
    .SDIN(n7420),
    .SDIN_t(n7420_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7421),
    .Q_t(n7421_t),
    .QN(n5638),
    .QN_t(n5638_t)
  );


  sdffs1
  \DFF_865/Q_reg 
  (
    .DIN(WX5946),
    .DIN_t(WX5946_t),
    .SDIN(n7419),
    .SDIN_t(n7419_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7420),
    .Q_t(n7420_t),
    .QN(n5643),
    .QN_t(n5643_t)
  );


  sdffs1
  \DFF_864/Q_reg 
  (
    .DIN(WX5944),
    .DIN_t(WX5944_t),
    .SDIN(n7418),
    .SDIN_t(n7418_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7419),
    .Q_t(n7419_t),
    .QN(n5648),
    .QN_t(n5648_t)
  );


  sdffs1
  \DFF_863/Q_reg 
  (
    .DIN(WX5942),
    .DIN_t(WX5942_t),
    .SDIN(n7417),
    .SDIN_t(n7417_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7418),
    .Q_t(n7418_t),
    .QN(n5508),
    .QN_t(n5508_t)
  );


  sdffs1
  \DFF_862/Q_reg 
  (
    .DIN(WX5940),
    .DIN_t(WX5940_t),
    .SDIN(n7416),
    .SDIN_t(n7416_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7417),
    .Q_t(n7417_t),
    .QN(n5512),
    .QN_t(n5512_t)
  );


  sdffs1
  \DFF_861/Q_reg 
  (
    .DIN(WX5938),
    .DIN_t(WX5938_t),
    .SDIN(n7415),
    .SDIN_t(n7415_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7416),
    .Q_t(n7416_t),
    .QN(n5516),
    .QN_t(n5516_t)
  );


  sdffs1
  \DFF_860/Q_reg 
  (
    .DIN(WX5936),
    .DIN_t(WX5936_t),
    .SDIN(n7414),
    .SDIN_t(n7414_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7415),
    .Q_t(n7415_t),
    .QN(n5520),
    .QN_t(n5520_t)
  );


  sdffs1
  \DFF_859/Q_reg 
  (
    .DIN(WX5934),
    .DIN_t(WX5934_t),
    .SDIN(n7413),
    .SDIN_t(n7413_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7414),
    .Q_t(n7414_t),
    .QN(n5524),
    .QN_t(n5524_t)
  );


  sdffs1
  \DFF_858/Q_reg 
  (
    .DIN(WX5932),
    .DIN_t(WX5932_t),
    .SDIN(n7412),
    .SDIN_t(n7412_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7413),
    .Q_t(n7413_t),
    .QN(n5528),
    .QN_t(n5528_t)
  );


  sdffs1
  \DFF_857/Q_reg 
  (
    .DIN(WX5930),
    .DIN_t(WX5930_t),
    .SDIN(n7411),
    .SDIN_t(n7411_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7412),
    .Q_t(n7412_t),
    .QN(n5532),
    .QN_t(n5532_t)
  );


  sdffs1
  \DFF_856/Q_reg 
  (
    .DIN(WX5928),
    .DIN_t(WX5928_t),
    .SDIN(n7410),
    .SDIN_t(n7410_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7411),
    .Q_t(n7411_t),
    .QN(n5536),
    .QN_t(n5536_t)
  );


  sdffs1
  \DFF_855/Q_reg 
  (
    .DIN(WX5926),
    .DIN_t(WX5926_t),
    .SDIN(n7409),
    .SDIN_t(n7409_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7410),
    .Q_t(n7410_t),
    .QN(n5540),
    .QN_t(n5540_t)
  );


  sdffs1
  \DFF_854/Q_reg 
  (
    .DIN(WX5924),
    .DIN_t(WX5924_t),
    .SDIN(n7408),
    .SDIN_t(n7408_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7409),
    .Q_t(n7409_t),
    .QN(n5544),
    .QN_t(n5544_t)
  );


  sdffs1
  \DFF_853/Q_reg 
  (
    .DIN(WX5922),
    .DIN_t(WX5922_t),
    .SDIN(n7407),
    .SDIN_t(n7407_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7408),
    .Q_t(n7408_t),
    .QN(n5548),
    .QN_t(n5548_t)
  );


  sdffs1
  \DFF_852/Q_reg 
  (
    .DIN(WX5920),
    .DIN_t(WX5920_t),
    .SDIN(n7406),
    .SDIN_t(n7406_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7407),
    .Q_t(n7407_t),
    .QN(n5552),
    .QN_t(n5552_t)
  );


  sdffs1
  \DFF_851/Q_reg 
  (
    .DIN(WX5918),
    .DIN_t(WX5918_t),
    .SDIN(n7405),
    .SDIN_t(n7405_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7406),
    .Q_t(n7406_t),
    .QN(n5556),
    .QN_t(n5556_t)
  );


  sdffs1
  \DFF_850/Q_reg 
  (
    .DIN(WX5916),
    .DIN_t(WX5916_t),
    .SDIN(n7404),
    .SDIN_t(n7404_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7405),
    .Q_t(n7405_t),
    .QN(n5560),
    .QN_t(n5560_t)
  );


  sdffs1
  \DFF_849/Q_reg 
  (
    .DIN(WX5914),
    .DIN_t(WX5914_t),
    .SDIN(n7403),
    .SDIN_t(n7403_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7404),
    .Q_t(n7404_t),
    .QN(n5564),
    .QN_t(n5564_t)
  );


  sdffs1
  \DFF_848/Q_reg 
  (
    .DIN(WX5912),
    .DIN_t(WX5912_t),
    .SDIN(n5572),
    .SDIN_t(n5572_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7403),
    .Q_t(n7403_t),
    .QN(n5568),
    .QN_t(n5568_t)
  );


  sdffs1
  \DFF_847/Q_reg 
  (
    .DIN(WX5910),
    .DIN_t(WX5910_t),
    .SDIN(n5577),
    .SDIN_t(n5577_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5572),
    .Q_t(n5572_t)
  );


  sdffs1
  \DFF_846/Q_reg 
  (
    .DIN(WX5908),
    .DIN_t(WX5908_t),
    .SDIN(n5582),
    .SDIN_t(n5582_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5577),
    .Q_t(n5577_t)
  );


  sdffs1
  \DFF_845/Q_reg 
  (
    .DIN(WX5906),
    .DIN_t(WX5906_t),
    .SDIN(n5587),
    .SDIN_t(n5587_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5582),
    .Q_t(n5582_t)
  );


  sdffs1
  \DFF_844/Q_reg 
  (
    .DIN(WX5904),
    .DIN_t(WX5904_t),
    .SDIN(n5592),
    .SDIN_t(n5592_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5587),
    .Q_t(n5587_t)
  );


  sdffs1
  \DFF_843/Q_reg 
  (
    .DIN(WX5902),
    .DIN_t(WX5902_t),
    .SDIN(n5597),
    .SDIN_t(n5597_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5592),
    .Q_t(n5592_t)
  );


  sdffs1
  \DFF_842/Q_reg 
  (
    .DIN(WX5900),
    .DIN_t(WX5900_t),
    .SDIN(n5602),
    .SDIN_t(n5602_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5597),
    .Q_t(n5597_t)
  );


  sdffs1
  \DFF_841/Q_reg 
  (
    .DIN(WX5898),
    .DIN_t(WX5898_t),
    .SDIN(n5607),
    .SDIN_t(n5607_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5602),
    .Q_t(n5602_t)
  );


  sdffs1
  \DFF_840/Q_reg 
  (
    .DIN(WX5896),
    .DIN_t(WX5896_t),
    .SDIN(n5612),
    .SDIN_t(n5612_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5607),
    .Q_t(n5607_t)
  );


  sdffs1
  \DFF_839/Q_reg 
  (
    .DIN(WX5894),
    .DIN_t(WX5894_t),
    .SDIN(n5617),
    .SDIN_t(n5617_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5612),
    .Q_t(n5612_t)
  );


  sdffs1
  \DFF_838/Q_reg 
  (
    .DIN(WX5892),
    .DIN_t(WX5892_t),
    .SDIN(n5622),
    .SDIN_t(n5622_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5617),
    .Q_t(n5617_t)
  );


  sdffs1
  \DFF_837/Q_reg 
  (
    .DIN(WX5890),
    .DIN_t(WX5890_t),
    .SDIN(n5627),
    .SDIN_t(n5627_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5622),
    .Q_t(n5622_t)
  );


  sdffs1
  \DFF_836/Q_reg 
  (
    .DIN(WX5888),
    .DIN_t(WX5888_t),
    .SDIN(n5632),
    .SDIN_t(n5632_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5627),
    .Q_t(n5627_t)
  );


  sdffs1
  \DFF_835/Q_reg 
  (
    .DIN(WX5886),
    .DIN_t(WX5886_t),
    .SDIN(n5637),
    .SDIN_t(n5637_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5632),
    .Q_t(n5632_t)
  );


  sdffs1
  \DFF_834/Q_reg 
  (
    .DIN(WX5884),
    .DIN_t(WX5884_t),
    .SDIN(n5642),
    .SDIN_t(n5642_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5637),
    .Q_t(n5637_t)
  );


  sdffs1
  \DFF_833/Q_reg 
  (
    .DIN(WX5882),
    .DIN_t(WX5882_t),
    .SDIN(n5647),
    .SDIN_t(n5647_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5642),
    .Q_t(n5642_t)
  );


  sdffs1
  \DFF_832/Q_reg 
  (
    .DIN(WX5880),
    .DIN_t(WX5880_t),
    .SDIN(n5507),
    .SDIN_t(n5507_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5647),
    .Q_t(n5647_t)
  );


  sdffs1
  \DFF_831/Q_reg 
  (
    .DIN(WX5878),
    .DIN_t(WX5878_t),
    .SDIN(n5511),
    .SDIN_t(n5511_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5507),
    .Q_t(n5507_t)
  );


  sdffs1
  \DFF_830/Q_reg 
  (
    .DIN(WX5876),
    .DIN_t(WX5876_t),
    .SDIN(n5515),
    .SDIN_t(n5515_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5511),
    .Q_t(n5511_t)
  );


  sdffs1
  \DFF_829/Q_reg 
  (
    .DIN(WX5874),
    .DIN_t(WX5874_t),
    .SDIN(n5519),
    .SDIN_t(n5519_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5515),
    .Q_t(n5515_t)
  );


  sdffs1
  \DFF_828/Q_reg 
  (
    .DIN(WX5872),
    .DIN_t(WX5872_t),
    .SDIN(n5523),
    .SDIN_t(n5523_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5519),
    .Q_t(n5519_t)
  );


  sdffs1
  \DFF_827/Q_reg 
  (
    .DIN(WX5870),
    .DIN_t(WX5870_t),
    .SDIN(n5527),
    .SDIN_t(n5527_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5523),
    .Q_t(n5523_t)
  );


  sdffs1
  \DFF_826/Q_reg 
  (
    .DIN(WX5868),
    .DIN_t(WX5868_t),
    .SDIN(n5531),
    .SDIN_t(n5531_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5527),
    .Q_t(n5527_t)
  );


  sdffs1
  \DFF_825/Q_reg 
  (
    .DIN(WX5866),
    .DIN_t(WX5866_t),
    .SDIN(n5535),
    .SDIN_t(n5535_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5531),
    .Q_t(n5531_t)
  );


  sdffs1
  \DFF_824/Q_reg 
  (
    .DIN(WX5864),
    .DIN_t(WX5864_t),
    .SDIN(n5539),
    .SDIN_t(n5539_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5535),
    .Q_t(n5535_t)
  );


  sdffs1
  \DFF_823/Q_reg 
  (
    .DIN(WX5862),
    .DIN_t(WX5862_t),
    .SDIN(n5543),
    .SDIN_t(n5543_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5539),
    .Q_t(n5539_t)
  );


  sdffs1
  \DFF_822/Q_reg 
  (
    .DIN(WX5860),
    .DIN_t(WX5860_t),
    .SDIN(n5547),
    .SDIN_t(n5547_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5543),
    .Q_t(n5543_t)
  );


  sdffs1
  \DFF_821/Q_reg 
  (
    .DIN(WX5858),
    .DIN_t(WX5858_t),
    .SDIN(n5551),
    .SDIN_t(n5551_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5547),
    .Q_t(n5547_t)
  );


  sdffs1
  \DFF_820/Q_reg 
  (
    .DIN(WX5856),
    .DIN_t(WX5856_t),
    .SDIN(n5555),
    .SDIN_t(n5555_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5551),
    .Q_t(n5551_t)
  );


  sdffs1
  \DFF_819/Q_reg 
  (
    .DIN(WX5854),
    .DIN_t(WX5854_t),
    .SDIN(n5559),
    .SDIN_t(n5559_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5555),
    .Q_t(n5555_t)
  );


  sdffs1
  \DFF_818/Q_reg 
  (
    .DIN(WX5852),
    .DIN_t(WX5852_t),
    .SDIN(n5563),
    .SDIN_t(n5563_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5559),
    .Q_t(n5559_t)
  );


  sdffs1
  \DFF_817/Q_reg 
  (
    .DIN(WX5850),
    .DIN_t(WX5850_t),
    .SDIN(n5567),
    .SDIN_t(n5567_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5563),
    .Q_t(n5563_t)
  );


  sdffs1
  \DFF_816/Q_reg 
  (
    .DIN(WX5848),
    .DIN_t(WX5848_t),
    .SDIN(n7402),
    .SDIN_t(n7402_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5567),
    .Q_t(n5567_t)
  );


  sdffs1
  \DFF_815/Q_reg 
  (
    .DIN(WX5846),
    .DIN_t(WX5846_t),
    .SDIN(n7401),
    .SDIN_t(n7401_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7402),
    .Q_t(n7402_t),
    .QN(n5571),
    .QN_t(n5571_t)
  );


  sdffs1
  \DFF_814/Q_reg 
  (
    .DIN(WX5844),
    .DIN_t(WX5844_t),
    .SDIN(n7400),
    .SDIN_t(n7400_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7401),
    .Q_t(n7401_t),
    .QN(n5576),
    .QN_t(n5576_t)
  );


  sdffs1
  \DFF_813/Q_reg 
  (
    .DIN(WX5842),
    .DIN_t(WX5842_t),
    .SDIN(n7399),
    .SDIN_t(n7399_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7400),
    .Q_t(n7400_t),
    .QN(n5581),
    .QN_t(n5581_t)
  );


  sdffs1
  \DFF_812/Q_reg 
  (
    .DIN(WX5840),
    .DIN_t(WX5840_t),
    .SDIN(n7398),
    .SDIN_t(n7398_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7399),
    .Q_t(n7399_t),
    .QN(n5586),
    .QN_t(n5586_t)
  );


  sdffs1
  \DFF_811/Q_reg 
  (
    .DIN(WX5838),
    .DIN_t(WX5838_t),
    .SDIN(n7397),
    .SDIN_t(n7397_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7398),
    .Q_t(n7398_t),
    .QN(n5591),
    .QN_t(n5591_t)
  );


  sdffs1
  \DFF_810/Q_reg 
  (
    .DIN(WX5836),
    .DIN_t(WX5836_t),
    .SDIN(n7396),
    .SDIN_t(n7396_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7397),
    .Q_t(n7397_t),
    .QN(n5596),
    .QN_t(n5596_t)
  );


  sdffs1
  \DFF_809/Q_reg 
  (
    .DIN(WX5834),
    .DIN_t(WX5834_t),
    .SDIN(n7395),
    .SDIN_t(n7395_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7396),
    .Q_t(n7396_t),
    .QN(n5601),
    .QN_t(n5601_t)
  );


  sdffs1
  \DFF_808/Q_reg 
  (
    .DIN(WX5832),
    .DIN_t(WX5832_t),
    .SDIN(n7394),
    .SDIN_t(n7394_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7395),
    .Q_t(n7395_t),
    .QN(n5606),
    .QN_t(n5606_t)
  );


  sdffs1
  \DFF_807/Q_reg 
  (
    .DIN(WX5830),
    .DIN_t(WX5830_t),
    .SDIN(n7393),
    .SDIN_t(n7393_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7394),
    .Q_t(n7394_t),
    .QN(n5611),
    .QN_t(n5611_t)
  );


  sdffs1
  \DFF_806/Q_reg 
  (
    .DIN(WX5828),
    .DIN_t(WX5828_t),
    .SDIN(n7392),
    .SDIN_t(n7392_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7393),
    .Q_t(n7393_t),
    .QN(n5616),
    .QN_t(n5616_t)
  );


  sdffs1
  \DFF_805/Q_reg 
  (
    .DIN(WX5826),
    .DIN_t(WX5826_t),
    .SDIN(n7391),
    .SDIN_t(n7391_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7392),
    .Q_t(n7392_t),
    .QN(n5621),
    .QN_t(n5621_t)
  );


  sdffs1
  \DFF_804/Q_reg 
  (
    .DIN(WX5824),
    .DIN_t(WX5824_t),
    .SDIN(n7390),
    .SDIN_t(n7390_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7391),
    .Q_t(n7391_t),
    .QN(n5626),
    .QN_t(n5626_t)
  );


  sdffs1
  \DFF_803/Q_reg 
  (
    .DIN(WX5822),
    .DIN_t(WX5822_t),
    .SDIN(n7389),
    .SDIN_t(n7389_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7390),
    .Q_t(n7390_t),
    .QN(n5631),
    .QN_t(n5631_t)
  );


  sdffs1
  \DFF_802/Q_reg 
  (
    .DIN(WX5820),
    .DIN_t(WX5820_t),
    .SDIN(n7388),
    .SDIN_t(n7388_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7389),
    .Q_t(n7389_t),
    .QN(n5636),
    .QN_t(n5636_t)
  );


  sdffs1
  \DFF_801/Q_reg 
  (
    .DIN(WX5818),
    .DIN_t(WX5818_t),
    .SDIN(n7387),
    .SDIN_t(n7387_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7388),
    .Q_t(n7388_t),
    .QN(n5641),
    .QN_t(n5641_t)
  );


  sdffs1
  \DFF_800/Q_reg 
  (
    .DIN(WX5816),
    .DIN_t(WX5816_t),
    .SDIN(n7386),
    .SDIN_t(n7386_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7387),
    .Q_t(n7387_t),
    .QN(n5646),
    .QN_t(n5646_t)
  );


  sdffs1
  \DFF_799/Q_reg 
  (
    .DIN(WX5718),
    .DIN_t(WX5718_t),
    .SDIN(n7385),
    .SDIN_t(n7385_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7386),
    .Q_t(n7386_t),
    .QN(n5476),
    .QN_t(n5476_t)
  );


  sdffs1
  \DFF_798/Q_reg 
  (
    .DIN(WX5716),
    .DIN_t(WX5716_t),
    .SDIN(n7384),
    .SDIN_t(n7384_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7385),
    .Q_t(n7385_t),
    .QN(n5477),
    .QN_t(n5477_t)
  );


  sdffs1
  \DFF_797/Q_reg 
  (
    .DIN(WX5714),
    .DIN_t(WX5714_t),
    .SDIN(n7383),
    .SDIN_t(n7383_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7384),
    .Q_t(n7384_t),
    .QN(n5478),
    .QN_t(n5478_t)
  );


  sdffs1
  \DFF_796/Q_reg 
  (
    .DIN(WX5712),
    .DIN_t(WX5712_t),
    .SDIN(n7382),
    .SDIN_t(n7382_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7383),
    .Q_t(n7383_t),
    .QN(n5479),
    .QN_t(n5479_t)
  );


  sdffs1
  \DFF_795/Q_reg 
  (
    .DIN(WX5710),
    .DIN_t(WX5710_t),
    .SDIN(n7381),
    .SDIN_t(n7381_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7382),
    .Q_t(n7382_t),
    .QN(n5480),
    .QN_t(n5480_t)
  );


  sdffs1
  \DFF_794/Q_reg 
  (
    .DIN(WX5708),
    .DIN_t(WX5708_t),
    .SDIN(n7380),
    .SDIN_t(n7380_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7381),
    .Q_t(n7381_t),
    .QN(n5481),
    .QN_t(n5481_t)
  );


  sdffs1
  \DFF_793/Q_reg 
  (
    .DIN(WX5706),
    .DIN_t(WX5706_t),
    .SDIN(n7379),
    .SDIN_t(n7379_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7380),
    .Q_t(n7380_t),
    .QN(n5482),
    .QN_t(n5482_t)
  );


  sdffs1
  \DFF_792/Q_reg 
  (
    .DIN(WX5704),
    .DIN_t(WX5704_t),
    .SDIN(n7378),
    .SDIN_t(n7378_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7379),
    .Q_t(n7379_t),
    .QN(n5483),
    .QN_t(n5483_t)
  );


  sdffs1
  \DFF_791/Q_reg 
  (
    .DIN(WX5702),
    .DIN_t(WX5702_t),
    .SDIN(n7377),
    .SDIN_t(n7377_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7378),
    .Q_t(n7378_t),
    .QN(n5484),
    .QN_t(n5484_t)
  );


  sdffs1
  \DFF_790/Q_reg 
  (
    .DIN(WX5700),
    .DIN_t(WX5700_t),
    .SDIN(n7376),
    .SDIN_t(n7376_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7377),
    .Q_t(n7377_t),
    .QN(n5485),
    .QN_t(n5485_t)
  );


  sdffs1
  \DFF_789/Q_reg 
  (
    .DIN(WX5698),
    .DIN_t(WX5698_t),
    .SDIN(n7375),
    .SDIN_t(n7375_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7376),
    .Q_t(n7376_t),
    .QN(n5486),
    .QN_t(n5486_t)
  );


  sdffs1
  \DFF_788/Q_reg 
  (
    .DIN(WX5696),
    .DIN_t(WX5696_t),
    .SDIN(n7374),
    .SDIN_t(n7374_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7375),
    .Q_t(n7375_t),
    .QN(n5487),
    .QN_t(n5487_t)
  );


  sdffs1
  \DFF_787/Q_reg 
  (
    .DIN(WX5694),
    .DIN_t(WX5694_t),
    .SDIN(n7373),
    .SDIN_t(n7373_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7374),
    .Q_t(n7374_t),
    .QN(n5488),
    .QN_t(n5488_t)
  );


  sdffs1
  \DFF_786/Q_reg 
  (
    .DIN(WX5692),
    .DIN_t(WX5692_t),
    .SDIN(n7372),
    .SDIN_t(n7372_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7373),
    .Q_t(n7373_t),
    .QN(n5489),
    .QN_t(n5489_t)
  );


  sdffs1
  \DFF_785/Q_reg 
  (
    .DIN(WX5690),
    .DIN_t(WX5690_t),
    .SDIN(n7371),
    .SDIN_t(n7371_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7372),
    .Q_t(n7372_t),
    .QN(n5490),
    .QN_t(n5490_t)
  );


  sdffs1
  \DFF_784/Q_reg 
  (
    .DIN(WX5688),
    .DIN_t(WX5688_t),
    .SDIN(n7370),
    .SDIN_t(n7370_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7371),
    .Q_t(n7371_t),
    .QN(n5491),
    .QN_t(n5491_t)
  );


  sdffs1
  \DFF_783/Q_reg 
  (
    .DIN(WX5686),
    .DIN_t(WX5686_t),
    .SDIN(n7369),
    .SDIN_t(n7369_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7370),
    .Q_t(n7370_t),
    .QN(n5492),
    .QN_t(n5492_t)
  );


  sdffs1
  \DFF_782/Q_reg 
  (
    .DIN(WX5684),
    .DIN_t(WX5684_t),
    .SDIN(n7368),
    .SDIN_t(n7368_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7369),
    .Q_t(n7369_t),
    .QN(n5493),
    .QN_t(n5493_t)
  );


  sdffs1
  \DFF_781/Q_reg 
  (
    .DIN(WX5682),
    .DIN_t(WX5682_t),
    .SDIN(n7367),
    .SDIN_t(n7367_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7368),
    .Q_t(n7368_t),
    .QN(n5494),
    .QN_t(n5494_t)
  );


  sdffs1
  \DFF_780/Q_reg 
  (
    .DIN(WX5680),
    .DIN_t(WX5680_t),
    .SDIN(n7366),
    .SDIN_t(n7366_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7367),
    .Q_t(n7367_t),
    .QN(n5495),
    .QN_t(n5495_t)
  );


  sdffs1
  \DFF_779/Q_reg 
  (
    .DIN(WX5678),
    .DIN_t(WX5678_t),
    .SDIN(n7365),
    .SDIN_t(n7365_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7366),
    .Q_t(n7366_t),
    .QN(n5496),
    .QN_t(n5496_t)
  );


  sdffs1
  \DFF_778/Q_reg 
  (
    .DIN(WX5676),
    .DIN_t(WX5676_t),
    .SDIN(n7364),
    .SDIN_t(n7364_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7365),
    .Q_t(n7365_t),
    .QN(n5497),
    .QN_t(n5497_t)
  );


  sdffs1
  \DFF_777/Q_reg 
  (
    .DIN(WX5674),
    .DIN_t(WX5674_t),
    .SDIN(n7363),
    .SDIN_t(n7363_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7364),
    .Q_t(n7364_t),
    .QN(n5498),
    .QN_t(n5498_t)
  );


  sdffs1
  \DFF_776/Q_reg 
  (
    .DIN(WX5672),
    .DIN_t(WX5672_t),
    .SDIN(n7362),
    .SDIN_t(n7362_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7363),
    .Q_t(n7363_t),
    .QN(n5499),
    .QN_t(n5499_t)
  );


  sdffs1
  \DFF_775/Q_reg 
  (
    .DIN(WX5670),
    .DIN_t(WX5670_t),
    .SDIN(n7361),
    .SDIN_t(n7361_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7362),
    .Q_t(n7362_t),
    .QN(n5500),
    .QN_t(n5500_t)
  );


  sdffs1
  \DFF_774/Q_reg 
  (
    .DIN(WX5668),
    .DIN_t(WX5668_t),
    .SDIN(n7360),
    .SDIN_t(n7360_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7361),
    .Q_t(n7361_t),
    .QN(n5501),
    .QN_t(n5501_t)
  );


  sdffs1
  \DFF_773/Q_reg 
  (
    .DIN(WX5666),
    .DIN_t(WX5666_t),
    .SDIN(n7359),
    .SDIN_t(n7359_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7360),
    .Q_t(n7360_t),
    .QN(n5502),
    .QN_t(n5502_t)
  );


  sdffs1
  \DFF_772/Q_reg 
  (
    .DIN(WX5664),
    .DIN_t(WX5664_t),
    .SDIN(n7358),
    .SDIN_t(n7358_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7359),
    .Q_t(n7359_t),
    .QN(n5503),
    .QN_t(n5503_t)
  );


  sdffs1
  \DFF_771/Q_reg 
  (
    .DIN(WX5662),
    .DIN_t(WX5662_t),
    .SDIN(n7357),
    .SDIN_t(n7357_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7358),
    .Q_t(n7358_t),
    .QN(n5504),
    .QN_t(n5504_t)
  );


  sdffs1
  \DFF_770/Q_reg 
  (
    .DIN(WX5660),
    .DIN_t(WX5660_t),
    .SDIN(n7356),
    .SDIN_t(n7356_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7357),
    .Q_t(n7357_t),
    .QN(n5505),
    .QN_t(n5505_t)
  );


  sdffs1
  \DFF_769/Q_reg 
  (
    .DIN(WX5658),
    .DIN_t(WX5658_t),
    .SDIN(n7355),
    .SDIN_t(n7355_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7356),
    .Q_t(n7356_t),
    .QN(n5506),
    .QN_t(n5506_t)
  );


  sdffs1
  \DFF_768/Q_reg 
  (
    .DIN(WX5656),
    .DIN_t(WX5656_t),
    .SDIN(CRC_OUT_6_31),
    .SDIN_t(CRC_OUT_6_31_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7355),
    .Q_t(n7355_t),
    .QN(n5475),
    .QN_t(n5475_t)
  );


  sdffs1
  \DFF_767/Q_reg 
  (
    .DIN(WX5205),
    .DIN_t(WX5205_t),
    .SDIN(CRC_OUT_6_30),
    .SDIN_t(CRC_OUT_6_30_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_31),
    .Q_t(CRC_OUT_6_31_t),
    .QN(n5650),
    .QN_t(n5650_t)
  );


  sdffs1
  \DFF_766/Q_reg 
  (
    .DIN(WX5203),
    .DIN_t(WX5203_t),
    .SDIN(CRC_OUT_6_29),
    .SDIN_t(CRC_OUT_6_29_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_30),
    .Q_t(CRC_OUT_6_30_t),
    .QN(n5645),
    .QN_t(n5645_t)
  );


  sdffs1
  \DFF_765/Q_reg 
  (
    .DIN(WX5201),
    .DIN_t(WX5201_t),
    .SDIN(CRC_OUT_6_28),
    .SDIN_t(CRC_OUT_6_28_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_29),
    .Q_t(CRC_OUT_6_29_t),
    .QN(n5640),
    .QN_t(n5640_t)
  );


  sdffs1
  \DFF_764/Q_reg 
  (
    .DIN(WX5199),
    .DIN_t(WX5199_t),
    .SDIN(CRC_OUT_6_27),
    .SDIN_t(CRC_OUT_6_27_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_28),
    .Q_t(CRC_OUT_6_28_t),
    .QN(n5635),
    .QN_t(n5635_t)
  );


  sdffs1
  \DFF_763/Q_reg 
  (
    .DIN(WX5197),
    .DIN_t(WX5197_t),
    .SDIN(CRC_OUT_6_26),
    .SDIN_t(CRC_OUT_6_26_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_27),
    .Q_t(CRC_OUT_6_27_t),
    .QN(n5630),
    .QN_t(n5630_t)
  );


  sdffs1
  \DFF_762/Q_reg 
  (
    .DIN(WX5195),
    .DIN_t(WX5195_t),
    .SDIN(CRC_OUT_6_25),
    .SDIN_t(CRC_OUT_6_25_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_26),
    .Q_t(CRC_OUT_6_26_t),
    .QN(n5625),
    .QN_t(n5625_t)
  );


  sdffs1
  \DFF_761/Q_reg 
  (
    .DIN(WX5193),
    .DIN_t(WX5193_t),
    .SDIN(CRC_OUT_6_24),
    .SDIN_t(CRC_OUT_6_24_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_25),
    .Q_t(CRC_OUT_6_25_t),
    .QN(n5620),
    .QN_t(n5620_t)
  );


  sdffs1
  \DFF_760/Q_reg 
  (
    .DIN(WX5191),
    .DIN_t(WX5191_t),
    .SDIN(CRC_OUT_6_23),
    .SDIN_t(CRC_OUT_6_23_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_24),
    .Q_t(CRC_OUT_6_24_t),
    .QN(n5615),
    .QN_t(n5615_t)
  );


  sdffs1
  \DFF_759/Q_reg 
  (
    .DIN(WX5189),
    .DIN_t(WX5189_t),
    .SDIN(CRC_OUT_6_22),
    .SDIN_t(CRC_OUT_6_22_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_23),
    .Q_t(CRC_OUT_6_23_t),
    .QN(n5610),
    .QN_t(n5610_t)
  );


  sdffs1
  \DFF_758/Q_reg 
  (
    .DIN(WX5187),
    .DIN_t(WX5187_t),
    .SDIN(CRC_OUT_6_21),
    .SDIN_t(CRC_OUT_6_21_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_22),
    .Q_t(CRC_OUT_6_22_t),
    .QN(n5605),
    .QN_t(n5605_t)
  );


  sdffs1
  \DFF_757/Q_reg 
  (
    .DIN(WX5185),
    .DIN_t(WX5185_t),
    .SDIN(CRC_OUT_6_20),
    .SDIN_t(CRC_OUT_6_20_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_21),
    .Q_t(CRC_OUT_6_21_t),
    .QN(n5600),
    .QN_t(n5600_t)
  );


  sdffs1
  \DFF_756/Q_reg 
  (
    .DIN(WX5183),
    .DIN_t(WX5183_t),
    .SDIN(CRC_OUT_6_19),
    .SDIN_t(CRC_OUT_6_19_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_20),
    .Q_t(CRC_OUT_6_20_t),
    .QN(n5595),
    .QN_t(n5595_t)
  );


  sdffs1
  \DFF_755/Q_reg 
  (
    .DIN(WX5181),
    .DIN_t(WX5181_t),
    .SDIN(CRC_OUT_6_18),
    .SDIN_t(CRC_OUT_6_18_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_19),
    .Q_t(CRC_OUT_6_19_t),
    .QN(n5590),
    .QN_t(n5590_t)
  );


  sdffs1
  \DFF_754/Q_reg 
  (
    .DIN(WX5179),
    .DIN_t(WX5179_t),
    .SDIN(CRC_OUT_6_17),
    .SDIN_t(CRC_OUT_6_17_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_18),
    .Q_t(CRC_OUT_6_18_t),
    .QN(n5585),
    .QN_t(n5585_t)
  );


  sdffs1
  \DFF_753/Q_reg 
  (
    .DIN(WX5177),
    .DIN_t(WX5177_t),
    .SDIN(CRC_OUT_6_16),
    .SDIN_t(CRC_OUT_6_16_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_17),
    .Q_t(CRC_OUT_6_17_t),
    .QN(n5580),
    .QN_t(n5580_t)
  );


  sdffs1
  \DFF_752/Q_reg 
  (
    .DIN(WX5175),
    .DIN_t(WX5175_t),
    .SDIN(CRC_OUT_6_15),
    .SDIN_t(CRC_OUT_6_15_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_16),
    .Q_t(CRC_OUT_6_16_t),
    .QN(n5575),
    .QN_t(n5575_t)
  );


  sdffs1
  \DFF_751/Q_reg 
  (
    .DIN(WX5173),
    .DIN_t(WX5173_t),
    .SDIN(CRC_OUT_6_14),
    .SDIN_t(CRC_OUT_6_14_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_15),
    .Q_t(CRC_OUT_6_15_t),
    .QN(n5570),
    .QN_t(n5570_t)
  );


  sdffs1
  \DFF_750/Q_reg 
  (
    .DIN(WX5171),
    .DIN_t(WX5171_t),
    .SDIN(CRC_OUT_6_13),
    .SDIN_t(CRC_OUT_6_13_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_14),
    .Q_t(CRC_OUT_6_14_t),
    .QN(n5566),
    .QN_t(n5566_t)
  );


  sdffs1
  \DFF_749/Q_reg 
  (
    .DIN(WX5169),
    .DIN_t(WX5169_t),
    .SDIN(CRC_OUT_6_12),
    .SDIN_t(CRC_OUT_6_12_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_13),
    .Q_t(CRC_OUT_6_13_t),
    .QN(n5562),
    .QN_t(n5562_t)
  );


  sdffs1
  \DFF_748/Q_reg 
  (
    .DIN(WX5167),
    .DIN_t(WX5167_t),
    .SDIN(CRC_OUT_6_11),
    .SDIN_t(CRC_OUT_6_11_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_12),
    .Q_t(CRC_OUT_6_12_t),
    .QN(n5558),
    .QN_t(n5558_t)
  );


  sdffs1
  \DFF_747/Q_reg 
  (
    .DIN(WX5165),
    .DIN_t(WX5165_t),
    .SDIN(CRC_OUT_6_10),
    .SDIN_t(CRC_OUT_6_10_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_11),
    .Q_t(CRC_OUT_6_11_t),
    .QN(n5554),
    .QN_t(n5554_t)
  );


  sdffs1
  \DFF_746/Q_reg 
  (
    .DIN(WX5163),
    .DIN_t(WX5163_t),
    .SDIN(CRC_OUT_6_9),
    .SDIN_t(CRC_OUT_6_9_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_10),
    .Q_t(CRC_OUT_6_10_t),
    .QN(n5550),
    .QN_t(n5550_t)
  );


  sdffs1
  \DFF_745/Q_reg 
  (
    .DIN(WX5161),
    .DIN_t(WX5161_t),
    .SDIN(CRC_OUT_6_8),
    .SDIN_t(CRC_OUT_6_8_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_9),
    .Q_t(CRC_OUT_6_9_t),
    .QN(n5546),
    .QN_t(n5546_t)
  );


  sdffs1
  \DFF_744/Q_reg 
  (
    .DIN(WX5159),
    .DIN_t(WX5159_t),
    .SDIN(CRC_OUT_6_7),
    .SDIN_t(CRC_OUT_6_7_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_8),
    .Q_t(CRC_OUT_6_8_t),
    .QN(n5542),
    .QN_t(n5542_t)
  );


  sdffs1
  \DFF_743/Q_reg 
  (
    .DIN(WX5157),
    .DIN_t(WX5157_t),
    .SDIN(CRC_OUT_6_6),
    .SDIN_t(CRC_OUT_6_6_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_7),
    .Q_t(CRC_OUT_6_7_t),
    .QN(n5538),
    .QN_t(n5538_t)
  );


  sdffs1
  \DFF_742/Q_reg 
  (
    .DIN(WX5155),
    .DIN_t(WX5155_t),
    .SDIN(CRC_OUT_6_5),
    .SDIN_t(CRC_OUT_6_5_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_6),
    .Q_t(CRC_OUT_6_6_t),
    .QN(n5534),
    .QN_t(n5534_t)
  );


  sdffs1
  \DFF_741/Q_reg 
  (
    .DIN(WX5153),
    .DIN_t(WX5153_t),
    .SDIN(CRC_OUT_6_4),
    .SDIN_t(CRC_OUT_6_4_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_5),
    .Q_t(CRC_OUT_6_5_t),
    .QN(n5530),
    .QN_t(n5530_t)
  );


  sdffs1
  \DFF_740/Q_reg 
  (
    .DIN(WX5151),
    .DIN_t(WX5151_t),
    .SDIN(CRC_OUT_6_3),
    .SDIN_t(CRC_OUT_6_3_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_4),
    .Q_t(CRC_OUT_6_4_t),
    .QN(n5526),
    .QN_t(n5526_t)
  );


  sdffs1
  \DFF_739/Q_reg 
  (
    .DIN(WX5149),
    .DIN_t(WX5149_t),
    .SDIN(CRC_OUT_6_2),
    .SDIN_t(CRC_OUT_6_2_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_3),
    .Q_t(CRC_OUT_6_3_t),
    .QN(n5522),
    .QN_t(n5522_t)
  );


  sdffs1
  \DFF_738/Q_reg 
  (
    .DIN(WX5147),
    .DIN_t(WX5147_t),
    .SDIN(CRC_OUT_6_1),
    .SDIN_t(CRC_OUT_6_1_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_2),
    .Q_t(CRC_OUT_6_2_t),
    .QN(n5518),
    .QN_t(n5518_t)
  );


  sdffs1
  \DFF_737/Q_reg 
  (
    .DIN(WX5145),
    .DIN_t(WX5145_t),
    .SDIN(CRC_OUT_6_0),
    .SDIN_t(CRC_OUT_6_0_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_1),
    .Q_t(CRC_OUT_6_1_t),
    .QN(n5514),
    .QN_t(n5514_t)
  );


  sdffs1
  \DFF_736/Q_reg 
  (
    .DIN(WX5143),
    .DIN_t(WX5143_t),
    .SDIN(n7354),
    .SDIN_t(n7354_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_6_0),
    .Q_t(CRC_OUT_6_0_t),
    .QN(n5510),
    .QN_t(n5510_t)
  );


  sdffs1
  \DFF_735/Q_reg 
  (
    .DIN(WX4777),
    .DIN_t(WX4777_t),
    .SDIN(n7353),
    .SDIN_t(n7353_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7354),
    .Q_t(n7354_t),
    .QN(n3269),
    .QN_t(n3269_t)
  );


  sdffs1
  \DFF_734/Q_reg 
  (
    .DIN(WX4775),
    .DIN_t(WX4775_t),
    .SDIN(n7352),
    .SDIN_t(n7352_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7353),
    .Q_t(n7353_t),
    .QN(n3270),
    .QN_t(n3270_t)
  );


  sdffs1
  \DFF_733/Q_reg 
  (
    .DIN(WX4773),
    .DIN_t(WX4773_t),
    .SDIN(n7351),
    .SDIN_t(n7351_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7352),
    .Q_t(n7352_t),
    .QN(n3271),
    .QN_t(n3271_t)
  );


  sdffs1
  \DFF_732/Q_reg 
  (
    .DIN(WX4771),
    .DIN_t(WX4771_t),
    .SDIN(n7350),
    .SDIN_t(n7350_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7351),
    .Q_t(n7351_t),
    .QN(n3272),
    .QN_t(n3272_t)
  );


  sdffs1
  \DFF_731/Q_reg 
  (
    .DIN(WX4769),
    .DIN_t(WX4769_t),
    .SDIN(n7349),
    .SDIN_t(n7349_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7350),
    .Q_t(n7350_t),
    .QN(n3273),
    .QN_t(n3273_t)
  );


  sdffs1
  \DFF_730/Q_reg 
  (
    .DIN(WX4767),
    .DIN_t(WX4767_t),
    .SDIN(n7348),
    .SDIN_t(n7348_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7349),
    .Q_t(n7349_t),
    .QN(n3274),
    .QN_t(n3274_t)
  );


  sdffs1
  \DFF_729/Q_reg 
  (
    .DIN(WX4765),
    .DIN_t(WX4765_t),
    .SDIN(n7347),
    .SDIN_t(n7347_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7348),
    .Q_t(n7348_t),
    .QN(n3275),
    .QN_t(n3275_t)
  );


  sdffs1
  \DFF_728/Q_reg 
  (
    .DIN(WX4763),
    .DIN_t(WX4763_t),
    .SDIN(n7346),
    .SDIN_t(n7346_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7347),
    .Q_t(n7347_t),
    .QN(n3276),
    .QN_t(n3276_t)
  );


  sdffs1
  \DFF_727/Q_reg 
  (
    .DIN(WX4761),
    .DIN_t(WX4761_t),
    .SDIN(n7345),
    .SDIN_t(n7345_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7346),
    .Q_t(n7346_t),
    .QN(n3277),
    .QN_t(n3277_t)
  );


  sdffs1
  \DFF_726/Q_reg 
  (
    .DIN(WX4759),
    .DIN_t(WX4759_t),
    .SDIN(n7344),
    .SDIN_t(n7344_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7345),
    .Q_t(n7345_t),
    .QN(n3278),
    .QN_t(n3278_t)
  );


  sdffs1
  \DFF_725/Q_reg 
  (
    .DIN(WX4757),
    .DIN_t(WX4757_t),
    .SDIN(n7343),
    .SDIN_t(n7343_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7344),
    .Q_t(n7344_t),
    .QN(n3279),
    .QN_t(n3279_t)
  );


  sdffs1
  \DFF_724/Q_reg 
  (
    .DIN(WX4755),
    .DIN_t(WX4755_t),
    .SDIN(n7342),
    .SDIN_t(n7342_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7343),
    .Q_t(n7343_t),
    .QN(n3280),
    .QN_t(n3280_t)
  );


  sdffs1
  \DFF_723/Q_reg 
  (
    .DIN(WX4753),
    .DIN_t(WX4753_t),
    .SDIN(n7341),
    .SDIN_t(n7341_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7342),
    .Q_t(n7342_t),
    .QN(n3281),
    .QN_t(n3281_t)
  );


  sdffs1
  \DFF_722/Q_reg 
  (
    .DIN(WX4751),
    .DIN_t(WX4751_t),
    .SDIN(n7340),
    .SDIN_t(n7340_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7341),
    .Q_t(n7341_t),
    .QN(n3282),
    .QN_t(n3282_t)
  );


  sdffs1
  \DFF_721/Q_reg 
  (
    .DIN(WX4749),
    .DIN_t(WX4749_t),
    .SDIN(n7339),
    .SDIN_t(n7339_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7340),
    .Q_t(n7340_t),
    .QN(n3283),
    .QN_t(n3283_t)
  );


  sdffs1
  \DFF_720/Q_reg 
  (
    .DIN(WX4747),
    .DIN_t(WX4747_t),
    .SDIN(n7338),
    .SDIN_t(n7338_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7339),
    .Q_t(n7339_t),
    .QN(n3284),
    .QN_t(n3284_t)
  );


  sdffs1
  \DFF_719/Q_reg 
  (
    .DIN(WX4745),
    .DIN_t(WX4745_t),
    .SDIN(n7337),
    .SDIN_t(n7337_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7338),
    .Q_t(n7338_t),
    .QN(n5750),
    .QN_t(n5750_t)
  );


  sdffs1
  \DFF_718/Q_reg 
  (
    .DIN(WX4743),
    .DIN_t(WX4743_t),
    .SDIN(n7336),
    .SDIN_t(n7336_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7337),
    .Q_t(n7337_t),
    .QN(n5755),
    .QN_t(n5755_t)
  );


  sdffs1
  \DFF_717/Q_reg 
  (
    .DIN(WX4741),
    .DIN_t(WX4741_t),
    .SDIN(n7335),
    .SDIN_t(n7335_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7336),
    .Q_t(n7336_t),
    .QN(n5760),
    .QN_t(n5760_t)
  );


  sdffs1
  \DFF_716/Q_reg 
  (
    .DIN(WX4739),
    .DIN_t(WX4739_t),
    .SDIN(n7334),
    .SDIN_t(n7334_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7335),
    .Q_t(n7335_t),
    .QN(n5765),
    .QN_t(n5765_t)
  );


  sdffs1
  \DFF_715/Q_reg 
  (
    .DIN(WX4737),
    .DIN_t(WX4737_t),
    .SDIN(n7333),
    .SDIN_t(n7333_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7334),
    .Q_t(n7334_t),
    .QN(n5770),
    .QN_t(n5770_t)
  );


  sdffs1
  \DFF_714/Q_reg 
  (
    .DIN(WX4735),
    .DIN_t(WX4735_t),
    .SDIN(n7332),
    .SDIN_t(n7332_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7333),
    .Q_t(n7333_t),
    .QN(n5775),
    .QN_t(n5775_t)
  );


  sdffs1
  \DFF_713/Q_reg 
  (
    .DIN(WX4733),
    .DIN_t(WX4733_t),
    .SDIN(n7331),
    .SDIN_t(n7331_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7332),
    .Q_t(n7332_t),
    .QN(n5780),
    .QN_t(n5780_t)
  );


  sdffs1
  \DFF_712/Q_reg 
  (
    .DIN(WX4731),
    .DIN_t(WX4731_t),
    .SDIN(n7330),
    .SDIN_t(n7330_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7331),
    .Q_t(n7331_t),
    .QN(n5785),
    .QN_t(n5785_t)
  );


  sdffs1
  \DFF_711/Q_reg 
  (
    .DIN(WX4729),
    .DIN_t(WX4729_t),
    .SDIN(n7329),
    .SDIN_t(n7329_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7330),
    .Q_t(n7330_t),
    .QN(n5790),
    .QN_t(n5790_t)
  );


  sdffs1
  \DFF_710/Q_reg 
  (
    .DIN(WX4727),
    .DIN_t(WX4727_t),
    .SDIN(n7328),
    .SDIN_t(n7328_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7329),
    .Q_t(n7329_t),
    .QN(n5795),
    .QN_t(n5795_t)
  );


  sdffs1
  \DFF_709/Q_reg 
  (
    .DIN(WX4725),
    .DIN_t(WX4725_t),
    .SDIN(n7327),
    .SDIN_t(n7327_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7328),
    .Q_t(n7328_t),
    .QN(n5800),
    .QN_t(n5800_t)
  );


  sdffs1
  \DFF_708/Q_reg 
  (
    .DIN(WX4723),
    .DIN_t(WX4723_t),
    .SDIN(n7326),
    .SDIN_t(n7326_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7327),
    .Q_t(n7327_t),
    .QN(n5805),
    .QN_t(n5805_t)
  );


  sdffs1
  \DFF_707/Q_reg 
  (
    .DIN(WX4721),
    .DIN_t(WX4721_t),
    .SDIN(n7325),
    .SDIN_t(n7325_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7326),
    .Q_t(n7326_t),
    .QN(n5810),
    .QN_t(n5810_t)
  );


  sdffs1
  \DFF_706/Q_reg 
  (
    .DIN(WX4719),
    .DIN_t(WX4719_t),
    .SDIN(n7324),
    .SDIN_t(n7324_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7325),
    .Q_t(n7325_t),
    .QN(n5815),
    .QN_t(n5815_t)
  );


  sdffs1
  \DFF_705/Q_reg 
  (
    .DIN(WX4717),
    .DIN_t(WX4717_t),
    .SDIN(n7323),
    .SDIN_t(n7323_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7324),
    .Q_t(n7324_t),
    .QN(n5820),
    .QN_t(n5820_t)
  );


  sdffs1
  \DFF_704/Q_reg 
  (
    .DIN(WX4715),
    .DIN_t(WX4715_t),
    .SDIN(n7322),
    .SDIN_t(n7322_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7323),
    .Q_t(n7323_t),
    .QN(n5825),
    .QN_t(n5825_t)
  );


  sdffs1
  \DFF_703/Q_reg 
  (
    .DIN(WX4713),
    .DIN_t(WX4713_t),
    .SDIN(n7321),
    .SDIN_t(n7321_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7322),
    .Q_t(n7322_t),
    .QN(n5685),
    .QN_t(n5685_t)
  );


  sdffs1
  \DFF_702/Q_reg 
  (
    .DIN(WX4711),
    .DIN_t(WX4711_t),
    .SDIN(n7320),
    .SDIN_t(n7320_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7321),
    .Q_t(n7321_t),
    .QN(n5689),
    .QN_t(n5689_t)
  );


  sdffs1
  \DFF_701/Q_reg 
  (
    .DIN(WX4709),
    .DIN_t(WX4709_t),
    .SDIN(n7319),
    .SDIN_t(n7319_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7320),
    .Q_t(n7320_t),
    .QN(n5693),
    .QN_t(n5693_t)
  );


  sdffs1
  \DFF_700/Q_reg 
  (
    .DIN(WX4707),
    .DIN_t(WX4707_t),
    .SDIN(n7318),
    .SDIN_t(n7318_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7319),
    .Q_t(n7319_t),
    .QN(n5697),
    .QN_t(n5697_t)
  );


  sdffs1
  \DFF_699/Q_reg 
  (
    .DIN(WX4705),
    .DIN_t(WX4705_t),
    .SDIN(n7317),
    .SDIN_t(n7317_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7318),
    .Q_t(n7318_t),
    .QN(n5701),
    .QN_t(n5701_t)
  );


  sdffs1
  \DFF_698/Q_reg 
  (
    .DIN(WX4703),
    .DIN_t(WX4703_t),
    .SDIN(n7316),
    .SDIN_t(n7316_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7317),
    .Q_t(n7317_t),
    .QN(n5705),
    .QN_t(n5705_t)
  );


  sdffs1
  \DFF_697/Q_reg 
  (
    .DIN(WX4701),
    .DIN_t(WX4701_t),
    .SDIN(n7315),
    .SDIN_t(n7315_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7316),
    .Q_t(n7316_t),
    .QN(n5709),
    .QN_t(n5709_t)
  );


  sdffs1
  \DFF_696/Q_reg 
  (
    .DIN(WX4699),
    .DIN_t(WX4699_t),
    .SDIN(n7314),
    .SDIN_t(n7314_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7315),
    .Q_t(n7315_t),
    .QN(n5713),
    .QN_t(n5713_t)
  );


  sdffs1
  \DFF_695/Q_reg 
  (
    .DIN(WX4697),
    .DIN_t(WX4697_t),
    .SDIN(n7313),
    .SDIN_t(n7313_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7314),
    .Q_t(n7314_t),
    .QN(n5717),
    .QN_t(n5717_t)
  );


  sdffs1
  \DFF_694/Q_reg 
  (
    .DIN(WX4695),
    .DIN_t(WX4695_t),
    .SDIN(n7312),
    .SDIN_t(n7312_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7313),
    .Q_t(n7313_t),
    .QN(n5721),
    .QN_t(n5721_t)
  );


  sdffs1
  \DFF_693/Q_reg 
  (
    .DIN(WX4693),
    .DIN_t(WX4693_t),
    .SDIN(n7311),
    .SDIN_t(n7311_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7312),
    .Q_t(n7312_t),
    .QN(n5725),
    .QN_t(n5725_t)
  );


  sdffs1
  \DFF_692/Q_reg 
  (
    .DIN(WX4691),
    .DIN_t(WX4691_t),
    .SDIN(n7310),
    .SDIN_t(n7310_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7311),
    .Q_t(n7311_t),
    .QN(n5729),
    .QN_t(n5729_t)
  );


  sdffs1
  \DFF_691/Q_reg 
  (
    .DIN(WX4689),
    .DIN_t(WX4689_t),
    .SDIN(n7309),
    .SDIN_t(n7309_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7310),
    .Q_t(n7310_t),
    .QN(n5733),
    .QN_t(n5733_t)
  );


  sdffs1
  \DFF_690/Q_reg 
  (
    .DIN(WX4687),
    .DIN_t(WX4687_t),
    .SDIN(n7308),
    .SDIN_t(n7308_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7309),
    .Q_t(n7309_t),
    .QN(n5737),
    .QN_t(n5737_t)
  );


  sdffs1
  \DFF_689/Q_reg 
  (
    .DIN(WX4685),
    .DIN_t(WX4685_t),
    .SDIN(n7307),
    .SDIN_t(n7307_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7308),
    .Q_t(n7308_t),
    .QN(n5741),
    .QN_t(n5741_t)
  );


  sdffs1
  \DFF_688/Q_reg 
  (
    .DIN(WX4683),
    .DIN_t(WX4683_t),
    .SDIN(n7306),
    .SDIN_t(n7306_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7307),
    .Q_t(n7307_t),
    .QN(n5745),
    .QN_t(n5745_t)
  );


  sdffs1
  \DFF_687/Q_reg 
  (
    .DIN(WX4681),
    .DIN_t(WX4681_t),
    .SDIN(n7305),
    .SDIN_t(n7305_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7306),
    .Q_t(n7306_t),
    .QN(n5749),
    .QN_t(n5749_t)
  );


  sdffs1
  \DFF_686/Q_reg 
  (
    .DIN(WX4679),
    .DIN_t(WX4679_t),
    .SDIN(n7304),
    .SDIN_t(n7304_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7305),
    .Q_t(n7305_t),
    .QN(n5754),
    .QN_t(n5754_t)
  );


  sdffs1
  \DFF_685/Q_reg 
  (
    .DIN(WX4677),
    .DIN_t(WX4677_t),
    .SDIN(n7303),
    .SDIN_t(n7303_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7304),
    .Q_t(n7304_t),
    .QN(n5759),
    .QN_t(n5759_t)
  );


  sdffs1
  \DFF_684/Q_reg 
  (
    .DIN(WX4675),
    .DIN_t(WX4675_t),
    .SDIN(n7302),
    .SDIN_t(n7302_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7303),
    .Q_t(n7303_t),
    .QN(n5764),
    .QN_t(n5764_t)
  );


  sdffs1
  \DFF_683/Q_reg 
  (
    .DIN(WX4673),
    .DIN_t(WX4673_t),
    .SDIN(n7301),
    .SDIN_t(n7301_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7302),
    .Q_t(n7302_t),
    .QN(n5769),
    .QN_t(n5769_t)
  );


  sdffs1
  \DFF_682/Q_reg 
  (
    .DIN(WX4671),
    .DIN_t(WX4671_t),
    .SDIN(n7300),
    .SDIN_t(n7300_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7301),
    .Q_t(n7301_t),
    .QN(n5774),
    .QN_t(n5774_t)
  );


  sdffs1
  \DFF_681/Q_reg 
  (
    .DIN(WX4669),
    .DIN_t(WX4669_t),
    .SDIN(n7299),
    .SDIN_t(n7299_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7300),
    .Q_t(n7300_t),
    .QN(n5779),
    .QN_t(n5779_t)
  );


  sdffs1
  \DFF_680/Q_reg 
  (
    .DIN(WX4667),
    .DIN_t(WX4667_t),
    .SDIN(n7298),
    .SDIN_t(n7298_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7299),
    .Q_t(n7299_t),
    .QN(n5784),
    .QN_t(n5784_t)
  );


  sdffs1
  \DFF_679/Q_reg 
  (
    .DIN(WX4665),
    .DIN_t(WX4665_t),
    .SDIN(n7297),
    .SDIN_t(n7297_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7298),
    .Q_t(n7298_t),
    .QN(n5789),
    .QN_t(n5789_t)
  );


  sdffs1
  \DFF_678/Q_reg 
  (
    .DIN(WX4663),
    .DIN_t(WX4663_t),
    .SDIN(n7296),
    .SDIN_t(n7296_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7297),
    .Q_t(n7297_t),
    .QN(n5794),
    .QN_t(n5794_t)
  );


  sdffs1
  \DFF_677/Q_reg 
  (
    .DIN(WX4661),
    .DIN_t(WX4661_t),
    .SDIN(n7295),
    .SDIN_t(n7295_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7296),
    .Q_t(n7296_t),
    .QN(n5799),
    .QN_t(n5799_t)
  );


  sdffs1
  \DFF_676/Q_reg 
  (
    .DIN(WX4659),
    .DIN_t(WX4659_t),
    .SDIN(n7294),
    .SDIN_t(n7294_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7295),
    .Q_t(n7295_t),
    .QN(n5804),
    .QN_t(n5804_t)
  );


  sdffs1
  \DFF_675/Q_reg 
  (
    .DIN(WX4657),
    .DIN_t(WX4657_t),
    .SDIN(n7293),
    .SDIN_t(n7293_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7294),
    .Q_t(n7294_t),
    .QN(n5809),
    .QN_t(n5809_t)
  );


  sdffs1
  \DFF_674/Q_reg 
  (
    .DIN(WX4655),
    .DIN_t(WX4655_t),
    .SDIN(n7292),
    .SDIN_t(n7292_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7293),
    .Q_t(n7293_t),
    .QN(n5814),
    .QN_t(n5814_t)
  );


  sdffs1
  \DFF_673/Q_reg 
  (
    .DIN(WX4653),
    .DIN_t(WX4653_t),
    .SDIN(n7291),
    .SDIN_t(n7291_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7292),
    .Q_t(n7292_t),
    .QN(n5819),
    .QN_t(n5819_t)
  );


  sdffs1
  \DFF_672/Q_reg 
  (
    .DIN(WX4651),
    .DIN_t(WX4651_t),
    .SDIN(n7290),
    .SDIN_t(n7290_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7291),
    .Q_t(n7291_t),
    .QN(n5824),
    .QN_t(n5824_t)
  );


  sdffs1
  \DFF_671/Q_reg 
  (
    .DIN(WX4649),
    .DIN_t(WX4649_t),
    .SDIN(n7289),
    .SDIN_t(n7289_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7290),
    .Q_t(n7290_t),
    .QN(n5684),
    .QN_t(n5684_t)
  );


  sdffs1
  \DFF_670/Q_reg 
  (
    .DIN(WX4647),
    .DIN_t(WX4647_t),
    .SDIN(n7288),
    .SDIN_t(n7288_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7289),
    .Q_t(n7289_t),
    .QN(n5688),
    .QN_t(n5688_t)
  );


  sdffs1
  \DFF_669/Q_reg 
  (
    .DIN(WX4645),
    .DIN_t(WX4645_t),
    .SDIN(n7287),
    .SDIN_t(n7287_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7288),
    .Q_t(n7288_t),
    .QN(n5692),
    .QN_t(n5692_t)
  );


  sdffs1
  \DFF_668/Q_reg 
  (
    .DIN(WX4643),
    .DIN_t(WX4643_t),
    .SDIN(n7286),
    .SDIN_t(n7286_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7287),
    .Q_t(n7287_t),
    .QN(n5696),
    .QN_t(n5696_t)
  );


  sdffs1
  \DFF_667/Q_reg 
  (
    .DIN(WX4641),
    .DIN_t(WX4641_t),
    .SDIN(n7285),
    .SDIN_t(n7285_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7286),
    .Q_t(n7286_t),
    .QN(n5700),
    .QN_t(n5700_t)
  );


  sdffs1
  \DFF_666/Q_reg 
  (
    .DIN(WX4639),
    .DIN_t(WX4639_t),
    .SDIN(n7284),
    .SDIN_t(n7284_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7285),
    .Q_t(n7285_t),
    .QN(n5704),
    .QN_t(n5704_t)
  );


  sdffs1
  \DFF_665/Q_reg 
  (
    .DIN(WX4637),
    .DIN_t(WX4637_t),
    .SDIN(n7283),
    .SDIN_t(n7283_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7284),
    .Q_t(n7284_t),
    .QN(n5708),
    .QN_t(n5708_t)
  );


  sdffs1
  \DFF_664/Q_reg 
  (
    .DIN(WX4635),
    .DIN_t(WX4635_t),
    .SDIN(n7282),
    .SDIN_t(n7282_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7283),
    .Q_t(n7283_t),
    .QN(n5712),
    .QN_t(n5712_t)
  );


  sdffs1
  \DFF_663/Q_reg 
  (
    .DIN(WX4633),
    .DIN_t(WX4633_t),
    .SDIN(n7281),
    .SDIN_t(n7281_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7282),
    .Q_t(n7282_t),
    .QN(n5716),
    .QN_t(n5716_t)
  );


  sdffs1
  \DFF_662/Q_reg 
  (
    .DIN(WX4631),
    .DIN_t(WX4631_t),
    .SDIN(n7280),
    .SDIN_t(n7280_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7281),
    .Q_t(n7281_t),
    .QN(n5720),
    .QN_t(n5720_t)
  );


  sdffs1
  \DFF_661/Q_reg 
  (
    .DIN(WX4629),
    .DIN_t(WX4629_t),
    .SDIN(n7279),
    .SDIN_t(n7279_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7280),
    .Q_t(n7280_t),
    .QN(n5724),
    .QN_t(n5724_t)
  );


  sdffs1
  \DFF_660/Q_reg 
  (
    .DIN(WX4627),
    .DIN_t(WX4627_t),
    .SDIN(n7278),
    .SDIN_t(n7278_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7279),
    .Q_t(n7279_t),
    .QN(n5728),
    .QN_t(n5728_t)
  );


  sdffs1
  \DFF_659/Q_reg 
  (
    .DIN(WX4625),
    .DIN_t(WX4625_t),
    .SDIN(n7277),
    .SDIN_t(n7277_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7278),
    .Q_t(n7278_t),
    .QN(n5732),
    .QN_t(n5732_t)
  );


  sdffs1
  \DFF_658/Q_reg 
  (
    .DIN(WX4623),
    .DIN_t(WX4623_t),
    .SDIN(n7276),
    .SDIN_t(n7276_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7277),
    .Q_t(n7277_t),
    .QN(n5736),
    .QN_t(n5736_t)
  );


  sdffs1
  \DFF_657/Q_reg 
  (
    .DIN(WX4621),
    .DIN_t(WX4621_t),
    .SDIN(n7275),
    .SDIN_t(n7275_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7276),
    .Q_t(n7276_t),
    .QN(n5740),
    .QN_t(n5740_t)
  );


  sdffs1
  \DFF_656/Q_reg 
  (
    .DIN(WX4619),
    .DIN_t(WX4619_t),
    .SDIN(n5748),
    .SDIN_t(n5748_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7275),
    .Q_t(n7275_t),
    .QN(n5744),
    .QN_t(n5744_t)
  );


  sdffs1
  \DFF_655/Q_reg 
  (
    .DIN(WX4617),
    .DIN_t(WX4617_t),
    .SDIN(n5753),
    .SDIN_t(n5753_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5748),
    .Q_t(n5748_t)
  );


  sdffs1
  \DFF_654/Q_reg 
  (
    .DIN(WX4615),
    .DIN_t(WX4615_t),
    .SDIN(n5758),
    .SDIN_t(n5758_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5753),
    .Q_t(n5753_t)
  );


  sdffs1
  \DFF_653/Q_reg 
  (
    .DIN(WX4613),
    .DIN_t(WX4613_t),
    .SDIN(n5763),
    .SDIN_t(n5763_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5758),
    .Q_t(n5758_t)
  );


  sdffs1
  \DFF_652/Q_reg 
  (
    .DIN(WX4611),
    .DIN_t(WX4611_t),
    .SDIN(n5768),
    .SDIN_t(n5768_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5763),
    .Q_t(n5763_t)
  );


  sdffs1
  \DFF_651/Q_reg 
  (
    .DIN(WX4609),
    .DIN_t(WX4609_t),
    .SDIN(n5773),
    .SDIN_t(n5773_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5768),
    .Q_t(n5768_t)
  );


  sdffs1
  \DFF_650/Q_reg 
  (
    .DIN(WX4607),
    .DIN_t(WX4607_t),
    .SDIN(n5778),
    .SDIN_t(n5778_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5773),
    .Q_t(n5773_t)
  );


  sdffs1
  \DFF_649/Q_reg 
  (
    .DIN(WX4605),
    .DIN_t(WX4605_t),
    .SDIN(n5783),
    .SDIN_t(n5783_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5778),
    .Q_t(n5778_t)
  );


  sdffs1
  \DFF_648/Q_reg 
  (
    .DIN(WX4603),
    .DIN_t(WX4603_t),
    .SDIN(n5788),
    .SDIN_t(n5788_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5783),
    .Q_t(n5783_t)
  );


  sdffs1
  \DFF_647/Q_reg 
  (
    .DIN(WX4601),
    .DIN_t(WX4601_t),
    .SDIN(n5793),
    .SDIN_t(n5793_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5788),
    .Q_t(n5788_t)
  );


  sdffs1
  \DFF_646/Q_reg 
  (
    .DIN(WX4599),
    .DIN_t(WX4599_t),
    .SDIN(n5798),
    .SDIN_t(n5798_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5793),
    .Q_t(n5793_t)
  );


  sdffs1
  \DFF_645/Q_reg 
  (
    .DIN(WX4597),
    .DIN_t(WX4597_t),
    .SDIN(n5803),
    .SDIN_t(n5803_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5798),
    .Q_t(n5798_t)
  );


  sdffs1
  \DFF_644/Q_reg 
  (
    .DIN(WX4595),
    .DIN_t(WX4595_t),
    .SDIN(n5808),
    .SDIN_t(n5808_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5803),
    .Q_t(n5803_t)
  );


  sdffs1
  \DFF_643/Q_reg 
  (
    .DIN(WX4593),
    .DIN_t(WX4593_t),
    .SDIN(n5813),
    .SDIN_t(n5813_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5808),
    .Q_t(n5808_t)
  );


  sdffs1
  \DFF_642/Q_reg 
  (
    .DIN(WX4591),
    .DIN_t(WX4591_t),
    .SDIN(n5818),
    .SDIN_t(n5818_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5813),
    .Q_t(n5813_t)
  );


  sdffs1
  \DFF_641/Q_reg 
  (
    .DIN(WX4589),
    .DIN_t(WX4589_t),
    .SDIN(n5823),
    .SDIN_t(n5823_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5818),
    .Q_t(n5818_t)
  );


  sdffs1
  \DFF_640/Q_reg 
  (
    .DIN(WX4587),
    .DIN_t(WX4587_t),
    .SDIN(n5683),
    .SDIN_t(n5683_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5823),
    .Q_t(n5823_t)
  );


  sdffs1
  \DFF_639/Q_reg 
  (
    .DIN(WX4585),
    .DIN_t(WX4585_t),
    .SDIN(n5687),
    .SDIN_t(n5687_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5683),
    .Q_t(n5683_t)
  );


  sdffs1
  \DFF_638/Q_reg 
  (
    .DIN(WX4583),
    .DIN_t(WX4583_t),
    .SDIN(n5691),
    .SDIN_t(n5691_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5687),
    .Q_t(n5687_t)
  );


  sdffs1
  \DFF_637/Q_reg 
  (
    .DIN(WX4581),
    .DIN_t(WX4581_t),
    .SDIN(n5695),
    .SDIN_t(n5695_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5691),
    .Q_t(n5691_t)
  );


  sdffs1
  \DFF_636/Q_reg 
  (
    .DIN(WX4579),
    .DIN_t(WX4579_t),
    .SDIN(n5699),
    .SDIN_t(n5699_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5695),
    .Q_t(n5695_t)
  );


  sdffs1
  \DFF_635/Q_reg 
  (
    .DIN(WX4577),
    .DIN_t(WX4577_t),
    .SDIN(n5703),
    .SDIN_t(n5703_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5699),
    .Q_t(n5699_t)
  );


  sdffs1
  \DFF_634/Q_reg 
  (
    .DIN(WX4575),
    .DIN_t(WX4575_t),
    .SDIN(n5707),
    .SDIN_t(n5707_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5703),
    .Q_t(n5703_t)
  );


  sdffs1
  \DFF_633/Q_reg 
  (
    .DIN(WX4573),
    .DIN_t(WX4573_t),
    .SDIN(n5711),
    .SDIN_t(n5711_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5707),
    .Q_t(n5707_t)
  );


  sdffs1
  \DFF_632/Q_reg 
  (
    .DIN(WX4571),
    .DIN_t(WX4571_t),
    .SDIN(n5715),
    .SDIN_t(n5715_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5711),
    .Q_t(n5711_t)
  );


  sdffs1
  \DFF_631/Q_reg 
  (
    .DIN(WX4569),
    .DIN_t(WX4569_t),
    .SDIN(n5719),
    .SDIN_t(n5719_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5715),
    .Q_t(n5715_t)
  );


  sdffs1
  \DFF_630/Q_reg 
  (
    .DIN(WX4567),
    .DIN_t(WX4567_t),
    .SDIN(n5723),
    .SDIN_t(n5723_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5719),
    .Q_t(n5719_t)
  );


  sdffs1
  \DFF_629/Q_reg 
  (
    .DIN(WX4565),
    .DIN_t(WX4565_t),
    .SDIN(n5727),
    .SDIN_t(n5727_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5723),
    .Q_t(n5723_t)
  );


  sdffs1
  \DFF_628/Q_reg 
  (
    .DIN(WX4563),
    .DIN_t(WX4563_t),
    .SDIN(n5731),
    .SDIN_t(n5731_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5727),
    .Q_t(n5727_t)
  );


  sdffs1
  \DFF_627/Q_reg 
  (
    .DIN(WX4561),
    .DIN_t(WX4561_t),
    .SDIN(n5735),
    .SDIN_t(n5735_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5731),
    .Q_t(n5731_t)
  );


  sdffs1
  \DFF_626/Q_reg 
  (
    .DIN(WX4559),
    .DIN_t(WX4559_t),
    .SDIN(n5739),
    .SDIN_t(n5739_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5735),
    .Q_t(n5735_t)
  );


  sdffs1
  \DFF_625/Q_reg 
  (
    .DIN(WX4557),
    .DIN_t(WX4557_t),
    .SDIN(n5743),
    .SDIN_t(n5743_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5739),
    .Q_t(n5739_t)
  );


  sdffs1
  \DFF_624/Q_reg 
  (
    .DIN(WX4555),
    .DIN_t(WX4555_t),
    .SDIN(n7274),
    .SDIN_t(n7274_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5743),
    .Q_t(n5743_t)
  );


  sdffs1
  \DFF_623/Q_reg 
  (
    .DIN(WX4553),
    .DIN_t(WX4553_t),
    .SDIN(n7273),
    .SDIN_t(n7273_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7274),
    .Q_t(n7274_t),
    .QN(n5747),
    .QN_t(n5747_t)
  );


  sdffs1
  \DFF_622/Q_reg 
  (
    .DIN(WX4551),
    .DIN_t(WX4551_t),
    .SDIN(n7272),
    .SDIN_t(n7272_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7273),
    .Q_t(n7273_t),
    .QN(n5752),
    .QN_t(n5752_t)
  );


  sdffs1
  \DFF_621/Q_reg 
  (
    .DIN(WX4549),
    .DIN_t(WX4549_t),
    .SDIN(n7271),
    .SDIN_t(n7271_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7272),
    .Q_t(n7272_t),
    .QN(n5757),
    .QN_t(n5757_t)
  );


  sdffs1
  \DFF_620/Q_reg 
  (
    .DIN(WX4547),
    .DIN_t(WX4547_t),
    .SDIN(n7270),
    .SDIN_t(n7270_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7271),
    .Q_t(n7271_t),
    .QN(n5762),
    .QN_t(n5762_t)
  );


  sdffs1
  \DFF_619/Q_reg 
  (
    .DIN(WX4545),
    .DIN_t(WX4545_t),
    .SDIN(n7269),
    .SDIN_t(n7269_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7270),
    .Q_t(n7270_t),
    .QN(n5767),
    .QN_t(n5767_t)
  );


  sdffs1
  \DFF_618/Q_reg 
  (
    .DIN(WX4543),
    .DIN_t(WX4543_t),
    .SDIN(n7268),
    .SDIN_t(n7268_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7269),
    .Q_t(n7269_t),
    .QN(n5772),
    .QN_t(n5772_t)
  );


  sdffs1
  \DFF_617/Q_reg 
  (
    .DIN(WX4541),
    .DIN_t(WX4541_t),
    .SDIN(n7267),
    .SDIN_t(n7267_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7268),
    .Q_t(n7268_t),
    .QN(n5777),
    .QN_t(n5777_t)
  );


  sdffs1
  \DFF_616/Q_reg 
  (
    .DIN(WX4539),
    .DIN_t(WX4539_t),
    .SDIN(n7266),
    .SDIN_t(n7266_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7267),
    .Q_t(n7267_t),
    .QN(n5782),
    .QN_t(n5782_t)
  );


  sdffs1
  \DFF_615/Q_reg 
  (
    .DIN(WX4537),
    .DIN_t(WX4537_t),
    .SDIN(n7265),
    .SDIN_t(n7265_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7266),
    .Q_t(n7266_t),
    .QN(n5787),
    .QN_t(n5787_t)
  );


  sdffs1
  \DFF_614/Q_reg 
  (
    .DIN(WX4535),
    .DIN_t(WX4535_t),
    .SDIN(n7264),
    .SDIN_t(n7264_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7265),
    .Q_t(n7265_t),
    .QN(n5792),
    .QN_t(n5792_t)
  );


  sdffs1
  \DFF_613/Q_reg 
  (
    .DIN(WX4533),
    .DIN_t(WX4533_t),
    .SDIN(n7263),
    .SDIN_t(n7263_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7264),
    .Q_t(n7264_t),
    .QN(n5797),
    .QN_t(n5797_t)
  );


  sdffs1
  \DFF_612/Q_reg 
  (
    .DIN(WX4531),
    .DIN_t(WX4531_t),
    .SDIN(n7262),
    .SDIN_t(n7262_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7263),
    .Q_t(n7263_t),
    .QN(n5802),
    .QN_t(n5802_t)
  );


  sdffs1
  \DFF_611/Q_reg 
  (
    .DIN(WX4529),
    .DIN_t(WX4529_t),
    .SDIN(n7261),
    .SDIN_t(n7261_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7262),
    .Q_t(n7262_t),
    .QN(n5807),
    .QN_t(n5807_t)
  );


  sdffs1
  \DFF_610/Q_reg 
  (
    .DIN(WX4527),
    .DIN_t(WX4527_t),
    .SDIN(n7260),
    .SDIN_t(n7260_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7261),
    .Q_t(n7261_t),
    .QN(n5812),
    .QN_t(n5812_t)
  );


  sdffs1
  \DFF_609/Q_reg 
  (
    .DIN(WX4525),
    .DIN_t(WX4525_t),
    .SDIN(n7259),
    .SDIN_t(n7259_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7260),
    .Q_t(n7260_t),
    .QN(n5817),
    .QN_t(n5817_t)
  );


  sdffs1
  \DFF_608/Q_reg 
  (
    .DIN(WX4523),
    .DIN_t(WX4523_t),
    .SDIN(n7258),
    .SDIN_t(n7258_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7259),
    .Q_t(n7259_t),
    .QN(n5822),
    .QN_t(n5822_t)
  );


  sdffs1
  \DFF_607/Q_reg 
  (
    .DIN(WX4425),
    .DIN_t(WX4425_t),
    .SDIN(n7257),
    .SDIN_t(n7257_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7258),
    .Q_t(n7258_t),
    .QN(n5652),
    .QN_t(n5652_t)
  );


  sdffs1
  \DFF_606/Q_reg 
  (
    .DIN(WX4423),
    .DIN_t(WX4423_t),
    .SDIN(n7256),
    .SDIN_t(n7256_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7257),
    .Q_t(n7257_t),
    .QN(n5653),
    .QN_t(n5653_t)
  );


  sdffs1
  \DFF_605/Q_reg 
  (
    .DIN(WX4421),
    .DIN_t(WX4421_t),
    .SDIN(n7255),
    .SDIN_t(n7255_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7256),
    .Q_t(n7256_t),
    .QN(n5654),
    .QN_t(n5654_t)
  );


  sdffs1
  \DFF_604/Q_reg 
  (
    .DIN(WX4419),
    .DIN_t(WX4419_t),
    .SDIN(n7254),
    .SDIN_t(n7254_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7255),
    .Q_t(n7255_t),
    .QN(n5655),
    .QN_t(n5655_t)
  );


  sdffs1
  \DFF_603/Q_reg 
  (
    .DIN(WX4417),
    .DIN_t(WX4417_t),
    .SDIN(n7253),
    .SDIN_t(n7253_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7254),
    .Q_t(n7254_t),
    .QN(n5656),
    .QN_t(n5656_t)
  );


  sdffs1
  \DFF_602/Q_reg 
  (
    .DIN(WX4415),
    .DIN_t(WX4415_t),
    .SDIN(n7252),
    .SDIN_t(n7252_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7253),
    .Q_t(n7253_t),
    .QN(n5657),
    .QN_t(n5657_t)
  );


  sdffs1
  \DFF_601/Q_reg 
  (
    .DIN(WX4413),
    .DIN_t(WX4413_t),
    .SDIN(n7251),
    .SDIN_t(n7251_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7252),
    .Q_t(n7252_t),
    .QN(n5658),
    .QN_t(n5658_t)
  );


  sdffs1
  \DFF_600/Q_reg 
  (
    .DIN(WX4411),
    .DIN_t(WX4411_t),
    .SDIN(n7250),
    .SDIN_t(n7250_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7251),
    .Q_t(n7251_t),
    .QN(n5659),
    .QN_t(n5659_t)
  );


  sdffs1
  \DFF_599/Q_reg 
  (
    .DIN(WX4409),
    .DIN_t(WX4409_t),
    .SDIN(n7249),
    .SDIN_t(n7249_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7250),
    .Q_t(n7250_t),
    .QN(n5660),
    .QN_t(n5660_t)
  );


  sdffs1
  \DFF_598/Q_reg 
  (
    .DIN(WX4407),
    .DIN_t(WX4407_t),
    .SDIN(n7248),
    .SDIN_t(n7248_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7249),
    .Q_t(n7249_t),
    .QN(n5661),
    .QN_t(n5661_t)
  );


  sdffs1
  \DFF_597/Q_reg 
  (
    .DIN(WX4405),
    .DIN_t(WX4405_t),
    .SDIN(n7247),
    .SDIN_t(n7247_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7248),
    .Q_t(n7248_t),
    .QN(n5662),
    .QN_t(n5662_t)
  );


  sdffs1
  \DFF_596/Q_reg 
  (
    .DIN(WX4403),
    .DIN_t(WX4403_t),
    .SDIN(n7246),
    .SDIN_t(n7246_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7247),
    .Q_t(n7247_t),
    .QN(n5663),
    .QN_t(n5663_t)
  );


  sdffs1
  \DFF_595/Q_reg 
  (
    .DIN(WX4401),
    .DIN_t(WX4401_t),
    .SDIN(n7245),
    .SDIN_t(n7245_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7246),
    .Q_t(n7246_t),
    .QN(n5664),
    .QN_t(n5664_t)
  );


  sdffs1
  \DFF_594/Q_reg 
  (
    .DIN(WX4399),
    .DIN_t(WX4399_t),
    .SDIN(n7244),
    .SDIN_t(n7244_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7245),
    .Q_t(n7245_t),
    .QN(n5665),
    .QN_t(n5665_t)
  );


  sdffs1
  \DFF_593/Q_reg 
  (
    .DIN(WX4397),
    .DIN_t(WX4397_t),
    .SDIN(n7243),
    .SDIN_t(n7243_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7244),
    .Q_t(n7244_t),
    .QN(n5666),
    .QN_t(n5666_t)
  );


  sdffs1
  \DFF_592/Q_reg 
  (
    .DIN(WX4395),
    .DIN_t(WX4395_t),
    .SDIN(n7242),
    .SDIN_t(n7242_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7243),
    .Q_t(n7243_t),
    .QN(n5667),
    .QN_t(n5667_t)
  );


  sdffs1
  \DFF_591/Q_reg 
  (
    .DIN(WX4393),
    .DIN_t(WX4393_t),
    .SDIN(n7241),
    .SDIN_t(n7241_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7242),
    .Q_t(n7242_t),
    .QN(n5668),
    .QN_t(n5668_t)
  );


  sdffs1
  \DFF_590/Q_reg 
  (
    .DIN(WX4391),
    .DIN_t(WX4391_t),
    .SDIN(n7240),
    .SDIN_t(n7240_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7241),
    .Q_t(n7241_t),
    .QN(n5669),
    .QN_t(n5669_t)
  );


  sdffs1
  \DFF_589/Q_reg 
  (
    .DIN(WX4389),
    .DIN_t(WX4389_t),
    .SDIN(n7239),
    .SDIN_t(n7239_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7240),
    .Q_t(n7240_t),
    .QN(n5670),
    .QN_t(n5670_t)
  );


  sdffs1
  \DFF_588/Q_reg 
  (
    .DIN(WX4387),
    .DIN_t(WX4387_t),
    .SDIN(n7238),
    .SDIN_t(n7238_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7239),
    .Q_t(n7239_t),
    .QN(n5671),
    .QN_t(n5671_t)
  );


  sdffs1
  \DFF_587/Q_reg 
  (
    .DIN(WX4385),
    .DIN_t(WX4385_t),
    .SDIN(n7237),
    .SDIN_t(n7237_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7238),
    .Q_t(n7238_t),
    .QN(n5672),
    .QN_t(n5672_t)
  );


  sdffs1
  \DFF_586/Q_reg 
  (
    .DIN(WX4383),
    .DIN_t(WX4383_t),
    .SDIN(n7236),
    .SDIN_t(n7236_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7237),
    .Q_t(n7237_t),
    .QN(n5673),
    .QN_t(n5673_t)
  );


  sdffs1
  \DFF_585/Q_reg 
  (
    .DIN(WX4381),
    .DIN_t(WX4381_t),
    .SDIN(n7235),
    .SDIN_t(n7235_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7236),
    .Q_t(n7236_t),
    .QN(n5674),
    .QN_t(n5674_t)
  );


  sdffs1
  \DFF_584/Q_reg 
  (
    .DIN(WX4379),
    .DIN_t(WX4379_t),
    .SDIN(n7234),
    .SDIN_t(n7234_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7235),
    .Q_t(n7235_t),
    .QN(n5675),
    .QN_t(n5675_t)
  );


  sdffs1
  \DFF_583/Q_reg 
  (
    .DIN(WX4377),
    .DIN_t(WX4377_t),
    .SDIN(n7233),
    .SDIN_t(n7233_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7234),
    .Q_t(n7234_t),
    .QN(n5676),
    .QN_t(n5676_t)
  );


  sdffs1
  \DFF_582/Q_reg 
  (
    .DIN(WX4375),
    .DIN_t(WX4375_t),
    .SDIN(n7232),
    .SDIN_t(n7232_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7233),
    .Q_t(n7233_t),
    .QN(n5677),
    .QN_t(n5677_t)
  );


  sdffs1
  \DFF_581/Q_reg 
  (
    .DIN(WX4373),
    .DIN_t(WX4373_t),
    .SDIN(n7231),
    .SDIN_t(n7231_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7232),
    .Q_t(n7232_t),
    .QN(n5678),
    .QN_t(n5678_t)
  );


  sdffs1
  \DFF_580/Q_reg 
  (
    .DIN(WX4371),
    .DIN_t(WX4371_t),
    .SDIN(n7230),
    .SDIN_t(n7230_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7231),
    .Q_t(n7231_t),
    .QN(n5679),
    .QN_t(n5679_t)
  );


  sdffs1
  \DFF_579/Q_reg 
  (
    .DIN(WX4369),
    .DIN_t(WX4369_t),
    .SDIN(n7229),
    .SDIN_t(n7229_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7230),
    .Q_t(n7230_t),
    .QN(n5680),
    .QN_t(n5680_t)
  );


  sdffs1
  \DFF_578/Q_reg 
  (
    .DIN(WX4367),
    .DIN_t(WX4367_t),
    .SDIN(n7228),
    .SDIN_t(n7228_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7229),
    .Q_t(n7229_t),
    .QN(n5681),
    .QN_t(n5681_t)
  );


  sdffs1
  \DFF_577/Q_reg 
  (
    .DIN(WX4365),
    .DIN_t(WX4365_t),
    .SDIN(n7227),
    .SDIN_t(n7227_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7228),
    .Q_t(n7228_t),
    .QN(n5682),
    .QN_t(n5682_t)
  );


  sdffs1
  \DFF_576/Q_reg 
  (
    .DIN(WX4363),
    .DIN_t(WX4363_t),
    .SDIN(CRC_OUT_7_31),
    .SDIN_t(CRC_OUT_7_31_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7227),
    .Q_t(n7227_t),
    .QN(n5651),
    .QN_t(n5651_t)
  );


  sdffs1
  \DFF_575/Q_reg 
  (
    .DIN(WX3912),
    .DIN_t(WX3912_t),
    .SDIN(CRC_OUT_7_30),
    .SDIN_t(CRC_OUT_7_30_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_31),
    .Q_t(CRC_OUT_7_31_t),
    .QN(n5826),
    .QN_t(n5826_t)
  );


  sdffs1
  \DFF_574/Q_reg 
  (
    .DIN(WX3910),
    .DIN_t(WX3910_t),
    .SDIN(CRC_OUT_7_29),
    .SDIN_t(CRC_OUT_7_29_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_30),
    .Q_t(CRC_OUT_7_30_t),
    .QN(n5821),
    .QN_t(n5821_t)
  );


  sdffs1
  \DFF_573/Q_reg 
  (
    .DIN(WX3908),
    .DIN_t(WX3908_t),
    .SDIN(CRC_OUT_7_28),
    .SDIN_t(CRC_OUT_7_28_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_29),
    .Q_t(CRC_OUT_7_29_t),
    .QN(n5816),
    .QN_t(n5816_t)
  );


  sdffs1
  \DFF_572/Q_reg 
  (
    .DIN(WX3906),
    .DIN_t(WX3906_t),
    .SDIN(CRC_OUT_7_27),
    .SDIN_t(CRC_OUT_7_27_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_28),
    .Q_t(CRC_OUT_7_28_t),
    .QN(n5811),
    .QN_t(n5811_t)
  );


  sdffs1
  \DFF_571/Q_reg 
  (
    .DIN(WX3904),
    .DIN_t(WX3904_t),
    .SDIN(CRC_OUT_7_26),
    .SDIN_t(CRC_OUT_7_26_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_27),
    .Q_t(CRC_OUT_7_27_t),
    .QN(n5806),
    .QN_t(n5806_t)
  );


  sdffs1
  \DFF_570/Q_reg 
  (
    .DIN(WX3902),
    .DIN_t(WX3902_t),
    .SDIN(CRC_OUT_7_25),
    .SDIN_t(CRC_OUT_7_25_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_26),
    .Q_t(CRC_OUT_7_26_t),
    .QN(n5801),
    .QN_t(n5801_t)
  );


  sdffs1
  \DFF_569/Q_reg 
  (
    .DIN(WX3900),
    .DIN_t(WX3900_t),
    .SDIN(CRC_OUT_7_24),
    .SDIN_t(CRC_OUT_7_24_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_25),
    .Q_t(CRC_OUT_7_25_t),
    .QN(n5796),
    .QN_t(n5796_t)
  );


  sdffs1
  \DFF_568/Q_reg 
  (
    .DIN(WX3898),
    .DIN_t(WX3898_t),
    .SDIN(CRC_OUT_7_23),
    .SDIN_t(CRC_OUT_7_23_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_24),
    .Q_t(CRC_OUT_7_24_t),
    .QN(n5791),
    .QN_t(n5791_t)
  );


  sdffs1
  \DFF_567/Q_reg 
  (
    .DIN(WX3896),
    .DIN_t(WX3896_t),
    .SDIN(CRC_OUT_7_22),
    .SDIN_t(CRC_OUT_7_22_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_23),
    .Q_t(CRC_OUT_7_23_t),
    .QN(n5786),
    .QN_t(n5786_t)
  );


  sdffs1
  \DFF_566/Q_reg 
  (
    .DIN(WX3894),
    .DIN_t(WX3894_t),
    .SDIN(CRC_OUT_7_21),
    .SDIN_t(CRC_OUT_7_21_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_22),
    .Q_t(CRC_OUT_7_22_t),
    .QN(n5781),
    .QN_t(n5781_t)
  );


  sdffs1
  \DFF_565/Q_reg 
  (
    .DIN(WX3892),
    .DIN_t(WX3892_t),
    .SDIN(CRC_OUT_7_20),
    .SDIN_t(CRC_OUT_7_20_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_21),
    .Q_t(CRC_OUT_7_21_t),
    .QN(n5776),
    .QN_t(n5776_t)
  );


  sdffs1
  \DFF_564/Q_reg 
  (
    .DIN(WX3890),
    .DIN_t(WX3890_t),
    .SDIN(CRC_OUT_7_19),
    .SDIN_t(CRC_OUT_7_19_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_20),
    .Q_t(CRC_OUT_7_20_t),
    .QN(n5771),
    .QN_t(n5771_t)
  );


  sdffs1
  \DFF_563/Q_reg 
  (
    .DIN(WX3888),
    .DIN_t(WX3888_t),
    .SDIN(CRC_OUT_7_18),
    .SDIN_t(CRC_OUT_7_18_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_19),
    .Q_t(CRC_OUT_7_19_t),
    .QN(n5766),
    .QN_t(n5766_t)
  );


  sdffs1
  \DFF_562/Q_reg 
  (
    .DIN(WX3886),
    .DIN_t(WX3886_t),
    .SDIN(CRC_OUT_7_17),
    .SDIN_t(CRC_OUT_7_17_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_18),
    .Q_t(CRC_OUT_7_18_t),
    .QN(n5761),
    .QN_t(n5761_t)
  );


  sdffs1
  \DFF_561/Q_reg 
  (
    .DIN(WX3884),
    .DIN_t(WX3884_t),
    .SDIN(CRC_OUT_7_16),
    .SDIN_t(CRC_OUT_7_16_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_17),
    .Q_t(CRC_OUT_7_17_t),
    .QN(n5756),
    .QN_t(n5756_t)
  );


  sdffs1
  \DFF_560/Q_reg 
  (
    .DIN(WX3882),
    .DIN_t(WX3882_t),
    .SDIN(CRC_OUT_7_15),
    .SDIN_t(CRC_OUT_7_15_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_16),
    .Q_t(CRC_OUT_7_16_t),
    .QN(n5751),
    .QN_t(n5751_t)
  );


  sdffs1
  \DFF_559/Q_reg 
  (
    .DIN(WX3880),
    .DIN_t(WX3880_t),
    .SDIN(CRC_OUT_7_14),
    .SDIN_t(CRC_OUT_7_14_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_15),
    .Q_t(CRC_OUT_7_15_t),
    .QN(n5746),
    .QN_t(n5746_t)
  );


  sdffs1
  \DFF_558/Q_reg 
  (
    .DIN(WX3878),
    .DIN_t(WX3878_t),
    .SDIN(CRC_OUT_7_13),
    .SDIN_t(CRC_OUT_7_13_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_14),
    .Q_t(CRC_OUT_7_14_t),
    .QN(n5742),
    .QN_t(n5742_t)
  );


  sdffs1
  \DFF_557/Q_reg 
  (
    .DIN(WX3876),
    .DIN_t(WX3876_t),
    .SDIN(CRC_OUT_7_12),
    .SDIN_t(CRC_OUT_7_12_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_13),
    .Q_t(CRC_OUT_7_13_t),
    .QN(n5738),
    .QN_t(n5738_t)
  );


  sdffs1
  \DFF_556/Q_reg 
  (
    .DIN(WX3874),
    .DIN_t(WX3874_t),
    .SDIN(CRC_OUT_7_11),
    .SDIN_t(CRC_OUT_7_11_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_12),
    .Q_t(CRC_OUT_7_12_t),
    .QN(n5734),
    .QN_t(n5734_t)
  );


  sdffs1
  \DFF_555/Q_reg 
  (
    .DIN(WX3872),
    .DIN_t(WX3872_t),
    .SDIN(CRC_OUT_7_10),
    .SDIN_t(CRC_OUT_7_10_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_11),
    .Q_t(CRC_OUT_7_11_t),
    .QN(n5730),
    .QN_t(n5730_t)
  );


  sdffs1
  \DFF_554/Q_reg 
  (
    .DIN(WX3870),
    .DIN_t(WX3870_t),
    .SDIN(CRC_OUT_7_9),
    .SDIN_t(CRC_OUT_7_9_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_10),
    .Q_t(CRC_OUT_7_10_t),
    .QN(n5726),
    .QN_t(n5726_t)
  );


  sdffs1
  \DFF_553/Q_reg 
  (
    .DIN(WX3868),
    .DIN_t(WX3868_t),
    .SDIN(CRC_OUT_7_8),
    .SDIN_t(CRC_OUT_7_8_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_9),
    .Q_t(CRC_OUT_7_9_t),
    .QN(n5722),
    .QN_t(n5722_t)
  );


  sdffs1
  \DFF_552/Q_reg 
  (
    .DIN(WX3866),
    .DIN_t(WX3866_t),
    .SDIN(CRC_OUT_7_7),
    .SDIN_t(CRC_OUT_7_7_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_8),
    .Q_t(CRC_OUT_7_8_t),
    .QN(n5718),
    .QN_t(n5718_t)
  );


  sdffs1
  \DFF_551/Q_reg 
  (
    .DIN(WX3864),
    .DIN_t(WX3864_t),
    .SDIN(CRC_OUT_7_6),
    .SDIN_t(CRC_OUT_7_6_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_7),
    .Q_t(CRC_OUT_7_7_t),
    .QN(n5714),
    .QN_t(n5714_t)
  );


  sdffs1
  \DFF_550/Q_reg 
  (
    .DIN(WX3862),
    .DIN_t(WX3862_t),
    .SDIN(CRC_OUT_7_5),
    .SDIN_t(CRC_OUT_7_5_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_6),
    .Q_t(CRC_OUT_7_6_t),
    .QN(n5710),
    .QN_t(n5710_t)
  );


  sdffs1
  \DFF_549/Q_reg 
  (
    .DIN(WX3860),
    .DIN_t(WX3860_t),
    .SDIN(CRC_OUT_7_4),
    .SDIN_t(CRC_OUT_7_4_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_5),
    .Q_t(CRC_OUT_7_5_t),
    .QN(n5706),
    .QN_t(n5706_t)
  );


  sdffs1
  \DFF_548/Q_reg 
  (
    .DIN(WX3858),
    .DIN_t(WX3858_t),
    .SDIN(CRC_OUT_7_3),
    .SDIN_t(CRC_OUT_7_3_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_4),
    .Q_t(CRC_OUT_7_4_t),
    .QN(n5702),
    .QN_t(n5702_t)
  );


  sdffs1
  \DFF_547/Q_reg 
  (
    .DIN(WX3856),
    .DIN_t(WX3856_t),
    .SDIN(CRC_OUT_7_2),
    .SDIN_t(CRC_OUT_7_2_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_3),
    .Q_t(CRC_OUT_7_3_t),
    .QN(n5698),
    .QN_t(n5698_t)
  );


  sdffs1
  \DFF_546/Q_reg 
  (
    .DIN(WX3854),
    .DIN_t(WX3854_t),
    .SDIN(CRC_OUT_7_1),
    .SDIN_t(CRC_OUT_7_1_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_2),
    .Q_t(CRC_OUT_7_2_t),
    .QN(n5694),
    .QN_t(n5694_t)
  );


  sdffs1
  \DFF_545/Q_reg 
  (
    .DIN(WX3852),
    .DIN_t(WX3852_t),
    .SDIN(CRC_OUT_7_0),
    .SDIN_t(CRC_OUT_7_0_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_1),
    .Q_t(CRC_OUT_7_1_t),
    .QN(n5690),
    .QN_t(n5690_t)
  );


  sdffs1
  \DFF_544/Q_reg 
  (
    .DIN(WX3850),
    .DIN_t(WX3850_t),
    .SDIN(n7226),
    .SDIN_t(n7226_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_7_0),
    .Q_t(CRC_OUT_7_0_t),
    .QN(n5686),
    .QN_t(n5686_t)
  );


  sdffs1
  \DFF_543/Q_reg 
  (
    .DIN(WX3484),
    .DIN_t(WX3484_t),
    .SDIN(n7225),
    .SDIN_t(n7225_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7226),
    .Q_t(n7226_t),
    .QN(n3285),
    .QN_t(n3285_t)
  );


  sdffs1
  \DFF_542/Q_reg 
  (
    .DIN(WX3482),
    .DIN_t(WX3482_t),
    .SDIN(n7224),
    .SDIN_t(n7224_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7225),
    .Q_t(n7225_t),
    .QN(n3287),
    .QN_t(n3287_t)
  );


  sdffs1
  \DFF_541/Q_reg 
  (
    .DIN(WX3480),
    .DIN_t(WX3480_t),
    .SDIN(n7223),
    .SDIN_t(n7223_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7224),
    .Q_t(n7224_t),
    .QN(n3289),
    .QN_t(n3289_t)
  );


  sdffs1
  \DFF_540/Q_reg 
  (
    .DIN(WX3478),
    .DIN_t(WX3478_t),
    .SDIN(n7222),
    .SDIN_t(n7222_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7223),
    .Q_t(n7223_t),
    .QN(n3291),
    .QN_t(n3291_t)
  );


  sdffs1
  \DFF_539/Q_reg 
  (
    .DIN(WX3476),
    .DIN_t(WX3476_t),
    .SDIN(n7221),
    .SDIN_t(n7221_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7222),
    .Q_t(n7222_t),
    .QN(n3293),
    .QN_t(n3293_t)
  );


  sdffs1
  \DFF_538/Q_reg 
  (
    .DIN(WX3474),
    .DIN_t(WX3474_t),
    .SDIN(n7220),
    .SDIN_t(n7220_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7221),
    .Q_t(n7221_t),
    .QN(n3295),
    .QN_t(n3295_t)
  );


  sdffs1
  \DFF_537/Q_reg 
  (
    .DIN(WX3472),
    .DIN_t(WX3472_t),
    .SDIN(n7219),
    .SDIN_t(n7219_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7220),
    .Q_t(n7220_t),
    .QN(n3297),
    .QN_t(n3297_t)
  );


  sdffs1
  \DFF_536/Q_reg 
  (
    .DIN(WX3470),
    .DIN_t(WX3470_t),
    .SDIN(n7218),
    .SDIN_t(n7218_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7219),
    .Q_t(n7219_t),
    .QN(n3299),
    .QN_t(n3299_t)
  );


  sdffs1
  \DFF_535/Q_reg 
  (
    .DIN(WX3468),
    .DIN_t(WX3468_t),
    .SDIN(n7217),
    .SDIN_t(n7217_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7218),
    .Q_t(n7218_t),
    .QN(n3301),
    .QN_t(n3301_t)
  );


  sdffs1
  \DFF_534/Q_reg 
  (
    .DIN(WX3466),
    .DIN_t(WX3466_t),
    .SDIN(n7216),
    .SDIN_t(n7216_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7217),
    .Q_t(n7217_t),
    .QN(n3303),
    .QN_t(n3303_t)
  );


  sdffs1
  \DFF_533/Q_reg 
  (
    .DIN(WX3464),
    .DIN_t(WX3464_t),
    .SDIN(n7215),
    .SDIN_t(n7215_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7216),
    .Q_t(n7216_t),
    .QN(n3305),
    .QN_t(n3305_t)
  );


  sdffs1
  \DFF_532/Q_reg 
  (
    .DIN(WX3462),
    .DIN_t(WX3462_t),
    .SDIN(n7214),
    .SDIN_t(n7214_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7215),
    .Q_t(n7215_t),
    .QN(n3307),
    .QN_t(n3307_t)
  );


  sdffs1
  \DFF_531/Q_reg 
  (
    .DIN(WX3460),
    .DIN_t(WX3460_t),
    .SDIN(n7213),
    .SDIN_t(n7213_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7214),
    .Q_t(n7214_t),
    .QN(n3309),
    .QN_t(n3309_t)
  );


  sdffs1
  \DFF_530/Q_reg 
  (
    .DIN(WX3458),
    .DIN_t(WX3458_t),
    .SDIN(n7212),
    .SDIN_t(n7212_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7213),
    .Q_t(n7213_t),
    .QN(n3311),
    .QN_t(n3311_t)
  );


  sdffs1
  \DFF_529/Q_reg 
  (
    .DIN(WX3456),
    .DIN_t(WX3456_t),
    .SDIN(n7211),
    .SDIN_t(n7211_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7212),
    .Q_t(n7212_t),
    .QN(n3313),
    .QN_t(n3313_t)
  );


  sdffs1
  \DFF_528/Q_reg 
  (
    .DIN(WX3454),
    .DIN_t(WX3454_t),
    .SDIN(n7210),
    .SDIN_t(n7210_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7211),
    .Q_t(n7211_t),
    .QN(n3315),
    .QN_t(n3315_t)
  );


  sdffs1
  \DFF_527/Q_reg 
  (
    .DIN(WX3452),
    .DIN_t(WX3452_t),
    .SDIN(n7209),
    .SDIN_t(n7209_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7210),
    .Q_t(n7210_t),
    .QN(n5974),
    .QN_t(n5974_t)
  );


  sdffs1
  \DFF_526/Q_reg 
  (
    .DIN(WX3450),
    .DIN_t(WX3450_t),
    .SDIN(n7208),
    .SDIN_t(n7208_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7209),
    .Q_t(n7209_t),
    .QN(n5983),
    .QN_t(n5983_t)
  );


  sdffs1
  \DFF_525/Q_reg 
  (
    .DIN(WX3448),
    .DIN_t(WX3448_t),
    .SDIN(n7207),
    .SDIN_t(n7207_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7208),
    .Q_t(n7208_t),
    .QN(n5992),
    .QN_t(n5992_t)
  );


  sdffs1
  \DFF_524/Q_reg 
  (
    .DIN(WX3446),
    .DIN_t(WX3446_t),
    .SDIN(n7206),
    .SDIN_t(n7206_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7207),
    .Q_t(n7207_t),
    .QN(n6001),
    .QN_t(n6001_t)
  );


  sdffs1
  \DFF_523/Q_reg 
  (
    .DIN(WX3444),
    .DIN_t(WX3444_t),
    .SDIN(n7205),
    .SDIN_t(n7205_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7206),
    .Q_t(n7206_t),
    .QN(n6010),
    .QN_t(n6010_t)
  );


  sdffs1
  \DFF_522/Q_reg 
  (
    .DIN(WX3442),
    .DIN_t(WX3442_t),
    .SDIN(n7204),
    .SDIN_t(n7204_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7205),
    .Q_t(n7205_t),
    .QN(n6019),
    .QN_t(n6019_t)
  );


  sdffs1
  \DFF_521/Q_reg 
  (
    .DIN(WX3440),
    .DIN_t(WX3440_t),
    .SDIN(n7203),
    .SDIN_t(n7203_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7204),
    .Q_t(n7204_t),
    .QN(n6028),
    .QN_t(n6028_t)
  );


  sdffs1
  \DFF_520/Q_reg 
  (
    .DIN(WX3438),
    .DIN_t(WX3438_t),
    .SDIN(n7202),
    .SDIN_t(n7202_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7203),
    .Q_t(n7203_t),
    .QN(n6037),
    .QN_t(n6037_t)
  );


  sdffs1
  \DFF_519/Q_reg 
  (
    .DIN(WX3436),
    .DIN_t(WX3436_t),
    .SDIN(n7201),
    .SDIN_t(n7201_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7202),
    .Q_t(n7202_t),
    .QN(n6046),
    .QN_t(n6046_t)
  );


  sdffs1
  \DFF_518/Q_reg 
  (
    .DIN(WX3434),
    .DIN_t(WX3434_t),
    .SDIN(n7200),
    .SDIN_t(n7200_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7201),
    .Q_t(n7201_t),
    .QN(n6055),
    .QN_t(n6055_t)
  );


  sdffs1
  \DFF_517/Q_reg 
  (
    .DIN(WX3432),
    .DIN_t(WX3432_t),
    .SDIN(n7199),
    .SDIN_t(n7199_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7200),
    .Q_t(n7200_t),
    .QN(n6064),
    .QN_t(n6064_t)
  );


  sdffs1
  \DFF_516/Q_reg 
  (
    .DIN(WX3430),
    .DIN_t(WX3430_t),
    .SDIN(n7198),
    .SDIN_t(n7198_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7199),
    .Q_t(n7199_t),
    .QN(n6073),
    .QN_t(n6073_t)
  );


  sdffs1
  \DFF_515/Q_reg 
  (
    .DIN(WX3428),
    .DIN_t(WX3428_t),
    .SDIN(n7197),
    .SDIN_t(n7197_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7198),
    .Q_t(n7198_t),
    .QN(n6082),
    .QN_t(n6082_t)
  );


  sdffs1
  \DFF_514/Q_reg 
  (
    .DIN(WX3426),
    .DIN_t(WX3426_t),
    .SDIN(n7196),
    .SDIN_t(n7196_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7197),
    .Q_t(n7197_t),
    .QN(n6091),
    .QN_t(n6091_t)
  );


  sdffs1
  \DFF_513/Q_reg 
  (
    .DIN(WX3424),
    .DIN_t(WX3424_t),
    .SDIN(n7195),
    .SDIN_t(n7195_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7196),
    .Q_t(n7196_t),
    .QN(n6100),
    .QN_t(n6100_t)
  );


  sdffs1
  \DFF_512/Q_reg 
  (
    .DIN(WX3422),
    .DIN_t(WX3422_t),
    .SDIN(n7194),
    .SDIN_t(n7194_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7195),
    .Q_t(n7195_t),
    .QN(n6109),
    .QN_t(n6109_t)
  );


  sdffs1
  \DFF_511/Q_reg 
  (
    .DIN(WX3420),
    .DIN_t(WX3420_t),
    .SDIN(n7193),
    .SDIN_t(n7193_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7194),
    .Q_t(n7194_t),
    .QN(n5861),
    .QN_t(n5861_t)
  );


  sdffs1
  \DFF_510/Q_reg 
  (
    .DIN(WX3418),
    .DIN_t(WX3418_t),
    .SDIN(n7192),
    .SDIN_t(n7192_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7193),
    .Q_t(n7193_t),
    .QN(n5868),
    .QN_t(n5868_t)
  );


  sdffs1
  \DFF_509/Q_reg 
  (
    .DIN(WX3416),
    .DIN_t(WX3416_t),
    .SDIN(n7191),
    .SDIN_t(n7191_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7192),
    .Q_t(n7192_t),
    .QN(n5875),
    .QN_t(n5875_t)
  );


  sdffs1
  \DFF_508/Q_reg 
  (
    .DIN(WX3414),
    .DIN_t(WX3414_t),
    .SDIN(n7190),
    .SDIN_t(n7190_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7191),
    .Q_t(n7191_t),
    .QN(n5882),
    .QN_t(n5882_t)
  );


  sdffs1
  \DFF_507/Q_reg 
  (
    .DIN(WX3412),
    .DIN_t(WX3412_t),
    .SDIN(n7189),
    .SDIN_t(n7189_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7190),
    .Q_t(n7190_t),
    .QN(n5889),
    .QN_t(n5889_t)
  );


  sdffs1
  \DFF_506/Q_reg 
  (
    .DIN(WX3410),
    .DIN_t(WX3410_t),
    .SDIN(n7188),
    .SDIN_t(n7188_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7189),
    .Q_t(n7189_t),
    .QN(n5896),
    .QN_t(n5896_t)
  );


  sdffs1
  \DFF_505/Q_reg 
  (
    .DIN(WX3408),
    .DIN_t(WX3408_t),
    .SDIN(n7187),
    .SDIN_t(n7187_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7188),
    .Q_t(n7188_t),
    .QN(n5903),
    .QN_t(n5903_t)
  );


  sdffs1
  \DFF_504/Q_reg 
  (
    .DIN(WX3406),
    .DIN_t(WX3406_t),
    .SDIN(n7186),
    .SDIN_t(n7186_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7187),
    .Q_t(n7187_t),
    .QN(n5910),
    .QN_t(n5910_t)
  );


  sdffs1
  \DFF_503/Q_reg 
  (
    .DIN(WX3404),
    .DIN_t(WX3404_t),
    .SDIN(n7185),
    .SDIN_t(n7185_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7186),
    .Q_t(n7186_t),
    .QN(n5917),
    .QN_t(n5917_t)
  );


  sdffs1
  \DFF_502/Q_reg 
  (
    .DIN(WX3402),
    .DIN_t(WX3402_t),
    .SDIN(n7184),
    .SDIN_t(n7184_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7185),
    .Q_t(n7185_t),
    .QN(n5924),
    .QN_t(n5924_t)
  );


  sdffs1
  \DFF_501/Q_reg 
  (
    .DIN(WX3400),
    .DIN_t(WX3400_t),
    .SDIN(n7183),
    .SDIN_t(n7183_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7184),
    .Q_t(n7184_t),
    .QN(n5931),
    .QN_t(n5931_t)
  );


  sdffs1
  \DFF_500/Q_reg 
  (
    .DIN(WX3398),
    .DIN_t(WX3398_t),
    .SDIN(n7182),
    .SDIN_t(n7182_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7183),
    .Q_t(n7183_t),
    .QN(n5938),
    .QN_t(n5938_t)
  );


  sdffs1
  \DFF_499/Q_reg 
  (
    .DIN(WX3396),
    .DIN_t(WX3396_t),
    .SDIN(n7181),
    .SDIN_t(n7181_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7182),
    .Q_t(n7182_t),
    .QN(n5945),
    .QN_t(n5945_t)
  );


  sdffs1
  \DFF_498/Q_reg 
  (
    .DIN(WX3394),
    .DIN_t(WX3394_t),
    .SDIN(n7180),
    .SDIN_t(n7180_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7181),
    .Q_t(n7181_t),
    .QN(n5952),
    .QN_t(n5952_t)
  );


  sdffs1
  \DFF_497/Q_reg 
  (
    .DIN(WX3392),
    .DIN_t(WX3392_t),
    .SDIN(n7179),
    .SDIN_t(n7179_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7180),
    .Q_t(n7180_t),
    .QN(n5959),
    .QN_t(n5959_t)
  );


  sdffs1
  \DFF_496/Q_reg 
  (
    .DIN(WX3390),
    .DIN_t(WX3390_t),
    .SDIN(n7178),
    .SDIN_t(n7178_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7179),
    .Q_t(n7179_t),
    .QN(n5966),
    .QN_t(n5966_t)
  );


  sdffs1
  \DFF_495/Q_reg 
  (
    .DIN(WX3388),
    .DIN_t(WX3388_t),
    .SDIN(n7177),
    .SDIN_t(n7177_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7178),
    .Q_t(n7178_t),
    .QN(n5973),
    .QN_t(n5973_t)
  );


  sdffs1
  \DFF_494/Q_reg 
  (
    .DIN(WX3386),
    .DIN_t(WX3386_t),
    .SDIN(n7176),
    .SDIN_t(n7176_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7177),
    .Q_t(n7177_t),
    .QN(n5982),
    .QN_t(n5982_t)
  );


  sdffs1
  \DFF_493/Q_reg 
  (
    .DIN(WX3384),
    .DIN_t(WX3384_t),
    .SDIN(n7175),
    .SDIN_t(n7175_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7176),
    .Q_t(n7176_t),
    .QN(n5991),
    .QN_t(n5991_t)
  );


  sdffs1
  \DFF_492/Q_reg 
  (
    .DIN(WX3382),
    .DIN_t(WX3382_t),
    .SDIN(n7174),
    .SDIN_t(n7174_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7175),
    .Q_t(n7175_t),
    .QN(n6000),
    .QN_t(n6000_t)
  );


  sdffs1
  \DFF_491/Q_reg 
  (
    .DIN(WX3380),
    .DIN_t(WX3380_t),
    .SDIN(n7173),
    .SDIN_t(n7173_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7174),
    .Q_t(n7174_t),
    .QN(n6009),
    .QN_t(n6009_t)
  );


  sdffs1
  \DFF_490/Q_reg 
  (
    .DIN(WX3378),
    .DIN_t(WX3378_t),
    .SDIN(n7172),
    .SDIN_t(n7172_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7173),
    .Q_t(n7173_t),
    .QN(n6018),
    .QN_t(n6018_t)
  );


  sdffs1
  \DFF_489/Q_reg 
  (
    .DIN(WX3376),
    .DIN_t(WX3376_t),
    .SDIN(n7171),
    .SDIN_t(n7171_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7172),
    .Q_t(n7172_t),
    .QN(n6027),
    .QN_t(n6027_t)
  );


  sdffs1
  \DFF_488/Q_reg 
  (
    .DIN(WX3374),
    .DIN_t(WX3374_t),
    .SDIN(n7170),
    .SDIN_t(n7170_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7171),
    .Q_t(n7171_t),
    .QN(n6036),
    .QN_t(n6036_t)
  );


  sdffs1
  \DFF_487/Q_reg 
  (
    .DIN(WX3372),
    .DIN_t(WX3372_t),
    .SDIN(n7169),
    .SDIN_t(n7169_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7170),
    .Q_t(n7170_t),
    .QN(n6045),
    .QN_t(n6045_t)
  );


  sdffs1
  \DFF_486/Q_reg 
  (
    .DIN(WX3370),
    .DIN_t(WX3370_t),
    .SDIN(n7168),
    .SDIN_t(n7168_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7169),
    .Q_t(n7169_t),
    .QN(n6054),
    .QN_t(n6054_t)
  );


  sdffs1
  \DFF_485/Q_reg 
  (
    .DIN(WX3368),
    .DIN_t(WX3368_t),
    .SDIN(n7167),
    .SDIN_t(n7167_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7168),
    .Q_t(n7168_t),
    .QN(n6063),
    .QN_t(n6063_t)
  );


  sdffs1
  \DFF_484/Q_reg 
  (
    .DIN(WX3366),
    .DIN_t(WX3366_t),
    .SDIN(n7166),
    .SDIN_t(n7166_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7167),
    .Q_t(n7167_t),
    .QN(n6072),
    .QN_t(n6072_t)
  );


  sdffs1
  \DFF_483/Q_reg 
  (
    .DIN(WX3364),
    .DIN_t(WX3364_t),
    .SDIN(n7165),
    .SDIN_t(n7165_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7166),
    .Q_t(n7166_t),
    .QN(n6081),
    .QN_t(n6081_t)
  );


  sdffs1
  \DFF_482/Q_reg 
  (
    .DIN(WX3362),
    .DIN_t(WX3362_t),
    .SDIN(n7164),
    .SDIN_t(n7164_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7165),
    .Q_t(n7165_t),
    .QN(n6090),
    .QN_t(n6090_t)
  );


  sdffs1
  \DFF_481/Q_reg 
  (
    .DIN(WX3360),
    .DIN_t(WX3360_t),
    .SDIN(n7163),
    .SDIN_t(n7163_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7164),
    .Q_t(n7164_t),
    .QN(n6099),
    .QN_t(n6099_t)
  );


  sdffs1
  \DFF_480/Q_reg 
  (
    .DIN(WX3358),
    .DIN_t(WX3358_t),
    .SDIN(n7162),
    .SDIN_t(n7162_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7163),
    .Q_t(n7163_t),
    .QN(n6108),
    .QN_t(n6108_t)
  );


  sdffs1
  \DFF_479/Q_reg 
  (
    .DIN(WX3356),
    .DIN_t(WX3356_t),
    .SDIN(n7161),
    .SDIN_t(n7161_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7162),
    .Q_t(n7162_t),
    .QN(n5860),
    .QN_t(n5860_t)
  );


  sdffs1
  \DFF_478/Q_reg 
  (
    .DIN(WX3354),
    .DIN_t(WX3354_t),
    .SDIN(n7160),
    .SDIN_t(n7160_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7161),
    .Q_t(n7161_t),
    .QN(n5867),
    .QN_t(n5867_t)
  );


  sdffs1
  \DFF_477/Q_reg 
  (
    .DIN(WX3352),
    .DIN_t(WX3352_t),
    .SDIN(n7159),
    .SDIN_t(n7159_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7160),
    .Q_t(n7160_t),
    .QN(n5874),
    .QN_t(n5874_t)
  );


  sdffs1
  \DFF_476/Q_reg 
  (
    .DIN(WX3350),
    .DIN_t(WX3350_t),
    .SDIN(n7158),
    .SDIN_t(n7158_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7159),
    .Q_t(n7159_t),
    .QN(n5881),
    .QN_t(n5881_t)
  );


  sdffs1
  \DFF_475/Q_reg 
  (
    .DIN(WX3348),
    .DIN_t(WX3348_t),
    .SDIN(n7157),
    .SDIN_t(n7157_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7158),
    .Q_t(n7158_t),
    .QN(n5888),
    .QN_t(n5888_t)
  );


  sdffs1
  \DFF_474/Q_reg 
  (
    .DIN(WX3346),
    .DIN_t(WX3346_t),
    .SDIN(n7156),
    .SDIN_t(n7156_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7157),
    .Q_t(n7157_t),
    .QN(n5895),
    .QN_t(n5895_t)
  );


  sdffs1
  \DFF_473/Q_reg 
  (
    .DIN(WX3344),
    .DIN_t(WX3344_t),
    .SDIN(n7155),
    .SDIN_t(n7155_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7156),
    .Q_t(n7156_t),
    .QN(n5902),
    .QN_t(n5902_t)
  );


  sdffs1
  \DFF_472/Q_reg 
  (
    .DIN(WX3342),
    .DIN_t(WX3342_t),
    .SDIN(n7154),
    .SDIN_t(n7154_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7155),
    .Q_t(n7155_t),
    .QN(n5909),
    .QN_t(n5909_t)
  );


  sdffs1
  \DFF_471/Q_reg 
  (
    .DIN(WX3340),
    .DIN_t(WX3340_t),
    .SDIN(n7153),
    .SDIN_t(n7153_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7154),
    .Q_t(n7154_t),
    .QN(n5916),
    .QN_t(n5916_t)
  );


  sdffs1
  \DFF_470/Q_reg 
  (
    .DIN(WX3338),
    .DIN_t(WX3338_t),
    .SDIN(n7152),
    .SDIN_t(n7152_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7153),
    .Q_t(n7153_t),
    .QN(n5923),
    .QN_t(n5923_t)
  );


  sdffs1
  \DFF_469/Q_reg 
  (
    .DIN(WX3336),
    .DIN_t(WX3336_t),
    .SDIN(n7151),
    .SDIN_t(n7151_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7152),
    .Q_t(n7152_t),
    .QN(n5930),
    .QN_t(n5930_t)
  );


  sdffs1
  \DFF_468/Q_reg 
  (
    .DIN(WX3334),
    .DIN_t(WX3334_t),
    .SDIN(n7150),
    .SDIN_t(n7150_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7151),
    .Q_t(n7151_t),
    .QN(n5937),
    .QN_t(n5937_t)
  );


  sdffs1
  \DFF_467/Q_reg 
  (
    .DIN(WX3332),
    .DIN_t(WX3332_t),
    .SDIN(n7149),
    .SDIN_t(n7149_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7150),
    .Q_t(n7150_t),
    .QN(n5944),
    .QN_t(n5944_t)
  );


  sdffs1
  \DFF_466/Q_reg 
  (
    .DIN(WX3330),
    .DIN_t(WX3330_t),
    .SDIN(n7148),
    .SDIN_t(n7148_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7149),
    .Q_t(n7149_t),
    .QN(n5951),
    .QN_t(n5951_t)
  );


  sdffs1
  \DFF_465/Q_reg 
  (
    .DIN(WX3328),
    .DIN_t(WX3328_t),
    .SDIN(n7147),
    .SDIN_t(n7147_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7148),
    .Q_t(n7148_t),
    .QN(n5958),
    .QN_t(n5958_t)
  );


  sdffs1
  \DFF_464/Q_reg 
  (
    .DIN(WX3326),
    .DIN_t(WX3326_t),
    .SDIN(n5972),
    .SDIN_t(n5972_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7147),
    .Q_t(n7147_t),
    .QN(n5965),
    .QN_t(n5965_t)
  );


  sdffs1
  \DFF_463/Q_reg 
  (
    .DIN(WX3324),
    .DIN_t(WX3324_t),
    .SDIN(n5981),
    .SDIN_t(n5981_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5972),
    .Q_t(n5972_t)
  );


  sdffs1
  \DFF_462/Q_reg 
  (
    .DIN(WX3322),
    .DIN_t(WX3322_t),
    .SDIN(n5990),
    .SDIN_t(n5990_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5981),
    .Q_t(n5981_t)
  );


  sdffs1
  \DFF_461/Q_reg 
  (
    .DIN(WX3320),
    .DIN_t(WX3320_t),
    .SDIN(n5999),
    .SDIN_t(n5999_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5990),
    .Q_t(n5990_t)
  );


  sdffs1
  \DFF_460/Q_reg 
  (
    .DIN(WX3318),
    .DIN_t(WX3318_t),
    .SDIN(n6008),
    .SDIN_t(n6008_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5999),
    .Q_t(n5999_t)
  );


  sdffs1
  \DFF_459/Q_reg 
  (
    .DIN(WX3316),
    .DIN_t(WX3316_t),
    .SDIN(n6017),
    .SDIN_t(n6017_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6008),
    .Q_t(n6008_t)
  );


  sdffs1
  \DFF_458/Q_reg 
  (
    .DIN(WX3314),
    .DIN_t(WX3314_t),
    .SDIN(n6026),
    .SDIN_t(n6026_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6017),
    .Q_t(n6017_t)
  );


  sdffs1
  \DFF_457/Q_reg 
  (
    .DIN(WX3312),
    .DIN_t(WX3312_t),
    .SDIN(n6035),
    .SDIN_t(n6035_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6026),
    .Q_t(n6026_t)
  );


  sdffs1
  \DFF_456/Q_reg 
  (
    .DIN(WX3310),
    .DIN_t(WX3310_t),
    .SDIN(n6044),
    .SDIN_t(n6044_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6035),
    .Q_t(n6035_t)
  );


  sdffs1
  \DFF_455/Q_reg 
  (
    .DIN(WX3308),
    .DIN_t(WX3308_t),
    .SDIN(n6053),
    .SDIN_t(n6053_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6044),
    .Q_t(n6044_t)
  );


  sdffs1
  \DFF_454/Q_reg 
  (
    .DIN(WX3306),
    .DIN_t(WX3306_t),
    .SDIN(n6062),
    .SDIN_t(n6062_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6053),
    .Q_t(n6053_t)
  );


  sdffs1
  \DFF_453/Q_reg 
  (
    .DIN(WX3304),
    .DIN_t(WX3304_t),
    .SDIN(n6071),
    .SDIN_t(n6071_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6062),
    .Q_t(n6062_t)
  );


  sdffs1
  \DFF_452/Q_reg 
  (
    .DIN(WX3302),
    .DIN_t(WX3302_t),
    .SDIN(n6080),
    .SDIN_t(n6080_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6071),
    .Q_t(n6071_t)
  );


  sdffs1
  \DFF_451/Q_reg 
  (
    .DIN(WX3300),
    .DIN_t(WX3300_t),
    .SDIN(n6089),
    .SDIN_t(n6089_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6080),
    .Q_t(n6080_t)
  );


  sdffs1
  \DFF_450/Q_reg 
  (
    .DIN(WX3298),
    .DIN_t(WX3298_t),
    .SDIN(n6098),
    .SDIN_t(n6098_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6089),
    .Q_t(n6089_t)
  );


  sdffs1
  \DFF_449/Q_reg 
  (
    .DIN(WX3296),
    .DIN_t(WX3296_t),
    .SDIN(n6107),
    .SDIN_t(n6107_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6098),
    .Q_t(n6098_t)
  );


  sdffs1
  \DFF_448/Q_reg 
  (
    .DIN(WX3294),
    .DIN_t(WX3294_t),
    .SDIN(n5859),
    .SDIN_t(n5859_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6107),
    .Q_t(n6107_t)
  );


  sdffs1
  \DFF_447/Q_reg 
  (
    .DIN(WX3292),
    .DIN_t(WX3292_t),
    .SDIN(n5866),
    .SDIN_t(n5866_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5859),
    .Q_t(n5859_t)
  );


  sdffs1
  \DFF_446/Q_reg 
  (
    .DIN(WX3290),
    .DIN_t(WX3290_t),
    .SDIN(n5873),
    .SDIN_t(n5873_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5866),
    .Q_t(n5866_t)
  );


  sdffs1
  \DFF_445/Q_reg 
  (
    .DIN(WX3288),
    .DIN_t(WX3288_t),
    .SDIN(n5880),
    .SDIN_t(n5880_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5873),
    .Q_t(n5873_t)
  );


  sdffs1
  \DFF_444/Q_reg 
  (
    .DIN(WX3286),
    .DIN_t(WX3286_t),
    .SDIN(n5887),
    .SDIN_t(n5887_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5880),
    .Q_t(n5880_t)
  );


  sdffs1
  \DFF_443/Q_reg 
  (
    .DIN(WX3284),
    .DIN_t(WX3284_t),
    .SDIN(n5894),
    .SDIN_t(n5894_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5887),
    .Q_t(n5887_t)
  );


  sdffs1
  \DFF_442/Q_reg 
  (
    .DIN(WX3282),
    .DIN_t(WX3282_t),
    .SDIN(n5901),
    .SDIN_t(n5901_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5894),
    .Q_t(n5894_t)
  );


  sdffs1
  \DFF_441/Q_reg 
  (
    .DIN(WX3280),
    .DIN_t(WX3280_t),
    .SDIN(n5908),
    .SDIN_t(n5908_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5901),
    .Q_t(n5901_t)
  );


  sdffs1
  \DFF_440/Q_reg 
  (
    .DIN(WX3278),
    .DIN_t(WX3278_t),
    .SDIN(n5915),
    .SDIN_t(n5915_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5908),
    .Q_t(n5908_t)
  );


  sdffs1
  \DFF_439/Q_reg 
  (
    .DIN(WX3276),
    .DIN_t(WX3276_t),
    .SDIN(n5922),
    .SDIN_t(n5922_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5915),
    .Q_t(n5915_t)
  );


  sdffs1
  \DFF_438/Q_reg 
  (
    .DIN(WX3274),
    .DIN_t(WX3274_t),
    .SDIN(n5929),
    .SDIN_t(n5929_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5922),
    .Q_t(n5922_t)
  );


  sdffs1
  \DFF_437/Q_reg 
  (
    .DIN(WX3272),
    .DIN_t(WX3272_t),
    .SDIN(n5936),
    .SDIN_t(n5936_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5929),
    .Q_t(n5929_t)
  );


  sdffs1
  \DFF_436/Q_reg 
  (
    .DIN(WX3270),
    .DIN_t(WX3270_t),
    .SDIN(n5943),
    .SDIN_t(n5943_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5936),
    .Q_t(n5936_t)
  );


  sdffs1
  \DFF_435/Q_reg 
  (
    .DIN(WX3268),
    .DIN_t(WX3268_t),
    .SDIN(n5950),
    .SDIN_t(n5950_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5943),
    .Q_t(n5943_t)
  );


  sdffs1
  \DFF_434/Q_reg 
  (
    .DIN(WX3266),
    .DIN_t(WX3266_t),
    .SDIN(n5957),
    .SDIN_t(n5957_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5950),
    .Q_t(n5950_t)
  );


  sdffs1
  \DFF_433/Q_reg 
  (
    .DIN(WX3264),
    .DIN_t(WX3264_t),
    .SDIN(n5964),
    .SDIN_t(n5964_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5957),
    .Q_t(n5957_t)
  );


  sdffs1
  \DFF_432/Q_reg 
  (
    .DIN(WX3262),
    .DIN_t(WX3262_t),
    .SDIN(n7146),
    .SDIN_t(n7146_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5964),
    .Q_t(n5964_t)
  );


  sdffs1
  \DFF_431/Q_reg 
  (
    .DIN(WX3260),
    .DIN_t(WX3260_t),
    .SDIN(n7145),
    .SDIN_t(n7145_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7146),
    .Q_t(n7146_t),
    .QN(n5971),
    .QN_t(n5971_t)
  );


  sdffs1
  \DFF_430/Q_reg 
  (
    .DIN(WX3258),
    .DIN_t(WX3258_t),
    .SDIN(n7144),
    .SDIN_t(n7144_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7145),
    .Q_t(n7145_t),
    .QN(n5980),
    .QN_t(n5980_t)
  );


  sdffs1
  \DFF_429/Q_reg 
  (
    .DIN(WX3256),
    .DIN_t(WX3256_t),
    .SDIN(n7143),
    .SDIN_t(n7143_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7144),
    .Q_t(n7144_t),
    .QN(n5989),
    .QN_t(n5989_t)
  );


  sdffs1
  \DFF_428/Q_reg 
  (
    .DIN(WX3254),
    .DIN_t(WX3254_t),
    .SDIN(n7142),
    .SDIN_t(n7142_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7143),
    .Q_t(n7143_t),
    .QN(n5998),
    .QN_t(n5998_t)
  );


  sdffs1
  \DFF_427/Q_reg 
  (
    .DIN(WX3252),
    .DIN_t(WX3252_t),
    .SDIN(n7141),
    .SDIN_t(n7141_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7142),
    .Q_t(n7142_t),
    .QN(n6007),
    .QN_t(n6007_t)
  );


  sdffs1
  \DFF_426/Q_reg 
  (
    .DIN(WX3250),
    .DIN_t(WX3250_t),
    .SDIN(n7140),
    .SDIN_t(n7140_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7141),
    .Q_t(n7141_t),
    .QN(n6016),
    .QN_t(n6016_t)
  );


  sdffs1
  \DFF_425/Q_reg 
  (
    .DIN(WX3248),
    .DIN_t(WX3248_t),
    .SDIN(n7139),
    .SDIN_t(n7139_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7140),
    .Q_t(n7140_t),
    .QN(n6025),
    .QN_t(n6025_t)
  );


  sdffs1
  \DFF_424/Q_reg 
  (
    .DIN(WX3246),
    .DIN_t(WX3246_t),
    .SDIN(n7138),
    .SDIN_t(n7138_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7139),
    .Q_t(n7139_t),
    .QN(n6034),
    .QN_t(n6034_t)
  );


  sdffs1
  \DFF_423/Q_reg 
  (
    .DIN(WX3244),
    .DIN_t(WX3244_t),
    .SDIN(n7137),
    .SDIN_t(n7137_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7138),
    .Q_t(n7138_t),
    .QN(n6043),
    .QN_t(n6043_t)
  );


  sdffs1
  \DFF_422/Q_reg 
  (
    .DIN(WX3242),
    .DIN_t(WX3242_t),
    .SDIN(n7136),
    .SDIN_t(n7136_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7137),
    .Q_t(n7137_t),
    .QN(n6052),
    .QN_t(n6052_t)
  );


  sdffs1
  \DFF_421/Q_reg 
  (
    .DIN(WX3240),
    .DIN_t(WX3240_t),
    .SDIN(n7135),
    .SDIN_t(n7135_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7136),
    .Q_t(n7136_t),
    .QN(n6061),
    .QN_t(n6061_t)
  );


  sdffs1
  \DFF_420/Q_reg 
  (
    .DIN(WX3238),
    .DIN_t(WX3238_t),
    .SDIN(n7134),
    .SDIN_t(n7134_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7135),
    .Q_t(n7135_t),
    .QN(n6070),
    .QN_t(n6070_t)
  );


  sdffs1
  \DFF_419/Q_reg 
  (
    .DIN(WX3236),
    .DIN_t(WX3236_t),
    .SDIN(n7133),
    .SDIN_t(n7133_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7134),
    .Q_t(n7134_t),
    .QN(n6079),
    .QN_t(n6079_t)
  );


  sdffs1
  \DFF_418/Q_reg 
  (
    .DIN(WX3234),
    .DIN_t(WX3234_t),
    .SDIN(n7132),
    .SDIN_t(n7132_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7133),
    .Q_t(n7133_t),
    .QN(n6088),
    .QN_t(n6088_t)
  );


  sdffs1
  \DFF_417/Q_reg 
  (
    .DIN(WX3232),
    .DIN_t(WX3232_t),
    .SDIN(n7131),
    .SDIN_t(n7131_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7132),
    .Q_t(n7132_t),
    .QN(n6097),
    .QN_t(n6097_t)
  );


  sdffs1
  \DFF_416/Q_reg 
  (
    .DIN(WX3230),
    .DIN_t(WX3230_t),
    .SDIN(n7130),
    .SDIN_t(n7130_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7131),
    .Q_t(n7131_t),
    .QN(n6106),
    .QN_t(n6106_t)
  );


  sdffs1
  \DFF_415/Q_reg 
  (
    .DIN(WX3132),
    .DIN_t(WX3132_t),
    .SDIN(n7129),
    .SDIN_t(n7129_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7130),
    .Q_t(n7130_t),
    .QN(n5828),
    .QN_t(n5828_t)
  );


  sdffs1
  \DFF_414/Q_reg 
  (
    .DIN(WX3130),
    .DIN_t(WX3130_t),
    .SDIN(n7128),
    .SDIN_t(n7128_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7129),
    .Q_t(n7129_t),
    .QN(n5829),
    .QN_t(n5829_t)
  );


  sdffs1
  \DFF_413/Q_reg 
  (
    .DIN(WX3128),
    .DIN_t(WX3128_t),
    .SDIN(n7127),
    .SDIN_t(n7127_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7128),
    .Q_t(n7128_t),
    .QN(n5830),
    .QN_t(n5830_t)
  );


  sdffs1
  \DFF_412/Q_reg 
  (
    .DIN(WX3126),
    .DIN_t(WX3126_t),
    .SDIN(n7126),
    .SDIN_t(n7126_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7127),
    .Q_t(n7127_t),
    .QN(n5831),
    .QN_t(n5831_t)
  );


  sdffs1
  \DFF_411/Q_reg 
  (
    .DIN(WX3124),
    .DIN_t(WX3124_t),
    .SDIN(n7125),
    .SDIN_t(n7125_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7126),
    .Q_t(n7126_t),
    .QN(n5832),
    .QN_t(n5832_t)
  );


  sdffs1
  \DFF_410/Q_reg 
  (
    .DIN(WX3122),
    .DIN_t(WX3122_t),
    .SDIN(n7124),
    .SDIN_t(n7124_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7125),
    .Q_t(n7125_t),
    .QN(n5833),
    .QN_t(n5833_t)
  );


  sdffs1
  \DFF_409/Q_reg 
  (
    .DIN(WX3120),
    .DIN_t(WX3120_t),
    .SDIN(n7123),
    .SDIN_t(n7123_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7124),
    .Q_t(n7124_t),
    .QN(n5834),
    .QN_t(n5834_t)
  );


  sdffs1
  \DFF_408/Q_reg 
  (
    .DIN(WX3118),
    .DIN_t(WX3118_t),
    .SDIN(n7122),
    .SDIN_t(n7122_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7123),
    .Q_t(n7123_t),
    .QN(n5835),
    .QN_t(n5835_t)
  );


  sdffs1
  \DFF_407/Q_reg 
  (
    .DIN(WX3116),
    .DIN_t(WX3116_t),
    .SDIN(n7121),
    .SDIN_t(n7121_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7122),
    .Q_t(n7122_t),
    .QN(n5836),
    .QN_t(n5836_t)
  );


  sdffs1
  \DFF_406/Q_reg 
  (
    .DIN(WX3114),
    .DIN_t(WX3114_t),
    .SDIN(n7120),
    .SDIN_t(n7120_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7121),
    .Q_t(n7121_t),
    .QN(n5837),
    .QN_t(n5837_t)
  );


  sdffs1
  \DFF_405/Q_reg 
  (
    .DIN(WX3112),
    .DIN_t(WX3112_t),
    .SDIN(n7119),
    .SDIN_t(n7119_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7120),
    .Q_t(n7120_t),
    .QN(n5838),
    .QN_t(n5838_t)
  );


  sdffs1
  \DFF_404/Q_reg 
  (
    .DIN(WX3110),
    .DIN_t(WX3110_t),
    .SDIN(n7118),
    .SDIN_t(n7118_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7119),
    .Q_t(n7119_t),
    .QN(n5839),
    .QN_t(n5839_t)
  );


  sdffs1
  \DFF_403/Q_reg 
  (
    .DIN(WX3108),
    .DIN_t(WX3108_t),
    .SDIN(n7117),
    .SDIN_t(n7117_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7118),
    .Q_t(n7118_t),
    .QN(n5840),
    .QN_t(n5840_t)
  );


  sdffs1
  \DFF_402/Q_reg 
  (
    .DIN(WX3106),
    .DIN_t(WX3106_t),
    .SDIN(n7116),
    .SDIN_t(n7116_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7117),
    .Q_t(n7117_t),
    .QN(n5841),
    .QN_t(n5841_t)
  );


  sdffs1
  \DFF_401/Q_reg 
  (
    .DIN(WX3104),
    .DIN_t(WX3104_t),
    .SDIN(n7115),
    .SDIN_t(n7115_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7116),
    .Q_t(n7116_t),
    .QN(n5842),
    .QN_t(n5842_t)
  );


  sdffs1
  \DFF_400/Q_reg 
  (
    .DIN(WX3102),
    .DIN_t(WX3102_t),
    .SDIN(n7114),
    .SDIN_t(n7114_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7115),
    .Q_t(n7115_t),
    .QN(n5843),
    .QN_t(n5843_t)
  );


  sdffs1
  \DFF_399/Q_reg 
  (
    .DIN(WX3100),
    .DIN_t(WX3100_t),
    .SDIN(n7113),
    .SDIN_t(n7113_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7114),
    .Q_t(n7114_t),
    .QN(n5844),
    .QN_t(n5844_t)
  );


  sdffs1
  \DFF_398/Q_reg 
  (
    .DIN(WX3098),
    .DIN_t(WX3098_t),
    .SDIN(n7112),
    .SDIN_t(n7112_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7113),
    .Q_t(n7113_t),
    .QN(n5845),
    .QN_t(n5845_t)
  );


  sdffs1
  \DFF_397/Q_reg 
  (
    .DIN(WX3096),
    .DIN_t(WX3096_t),
    .SDIN(n7111),
    .SDIN_t(n7111_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7112),
    .Q_t(n7112_t),
    .QN(n5846),
    .QN_t(n5846_t)
  );


  sdffs1
  \DFF_396/Q_reg 
  (
    .DIN(WX3094),
    .DIN_t(WX3094_t),
    .SDIN(n7110),
    .SDIN_t(n7110_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7111),
    .Q_t(n7111_t),
    .QN(n5847),
    .QN_t(n5847_t)
  );


  sdffs1
  \DFF_395/Q_reg 
  (
    .DIN(WX3092),
    .DIN_t(WX3092_t),
    .SDIN(n7109),
    .SDIN_t(n7109_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7110),
    .Q_t(n7110_t),
    .QN(n5848),
    .QN_t(n5848_t)
  );


  sdffs1
  \DFF_394/Q_reg 
  (
    .DIN(WX3090),
    .DIN_t(WX3090_t),
    .SDIN(n7108),
    .SDIN_t(n7108_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7109),
    .Q_t(n7109_t),
    .QN(n5849),
    .QN_t(n5849_t)
  );


  sdffs1
  \DFF_393/Q_reg 
  (
    .DIN(WX3088),
    .DIN_t(WX3088_t),
    .SDIN(n7107),
    .SDIN_t(n7107_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7108),
    .Q_t(n7108_t),
    .QN(n5850),
    .QN_t(n5850_t)
  );


  sdffs1
  \DFF_392/Q_reg 
  (
    .DIN(WX3086),
    .DIN_t(WX3086_t),
    .SDIN(n7106),
    .SDIN_t(n7106_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7107),
    .Q_t(n7107_t),
    .QN(n5851),
    .QN_t(n5851_t)
  );


  sdffs1
  \DFF_391/Q_reg 
  (
    .DIN(WX3084),
    .DIN_t(WX3084_t),
    .SDIN(n7105),
    .SDIN_t(n7105_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7106),
    .Q_t(n7106_t),
    .QN(n5852),
    .QN_t(n5852_t)
  );


  sdffs1
  \DFF_390/Q_reg 
  (
    .DIN(WX3082),
    .DIN_t(WX3082_t),
    .SDIN(n7104),
    .SDIN_t(n7104_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7105),
    .Q_t(n7105_t),
    .QN(n5853),
    .QN_t(n5853_t)
  );


  sdffs1
  \DFF_389/Q_reg 
  (
    .DIN(WX3080),
    .DIN_t(WX3080_t),
    .SDIN(n7103),
    .SDIN_t(n7103_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7104),
    .Q_t(n7104_t),
    .QN(n5854),
    .QN_t(n5854_t)
  );


  sdffs1
  \DFF_388/Q_reg 
  (
    .DIN(WX3078),
    .DIN_t(WX3078_t),
    .SDIN(n7102),
    .SDIN_t(n7102_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7103),
    .Q_t(n7103_t),
    .QN(n5855),
    .QN_t(n5855_t)
  );


  sdffs1
  \DFF_387/Q_reg 
  (
    .DIN(WX3076),
    .DIN_t(WX3076_t),
    .SDIN(n7101),
    .SDIN_t(n7101_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7102),
    .Q_t(n7102_t),
    .QN(n5856),
    .QN_t(n5856_t)
  );


  sdffs1
  \DFF_386/Q_reg 
  (
    .DIN(WX3074),
    .DIN_t(WX3074_t),
    .SDIN(n7100),
    .SDIN_t(n7100_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7101),
    .Q_t(n7101_t),
    .QN(n5857),
    .QN_t(n5857_t)
  );


  sdffs1
  \DFF_385/Q_reg 
  (
    .DIN(WX3072),
    .DIN_t(WX3072_t),
    .SDIN(n7099),
    .SDIN_t(n7099_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7100),
    .Q_t(n7100_t),
    .QN(n5858),
    .QN_t(n5858_t)
  );


  sdffs1
  \DFF_384/Q_reg 
  (
    .DIN(WX3070),
    .DIN_t(WX3070_t),
    .SDIN(CRC_OUT_8_31),
    .SDIN_t(CRC_OUT_8_31_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7099),
    .Q_t(n7099_t),
    .QN(n5827),
    .QN_t(n5827_t)
  );


  sdffs1
  \DFF_383/Q_reg 
  (
    .DIN(WX2619),
    .DIN_t(WX2619_t),
    .SDIN(CRC_OUT_8_30),
    .SDIN_t(CRC_OUT_8_30_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_31),
    .Q_t(CRC_OUT_8_31_t),
    .QN(n6114),
    .QN_t(n6114_t)
  );


  sdffs1
  \DFF_382/Q_reg 
  (
    .DIN(WX2617),
    .DIN_t(WX2617_t),
    .SDIN(CRC_OUT_8_29),
    .SDIN_t(CRC_OUT_8_29_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_30),
    .Q_t(CRC_OUT_8_30_t),
    .QN(n6105),
    .QN_t(n6105_t)
  );


  sdffs1
  \DFF_381/Q_reg 
  (
    .DIN(WX2615),
    .DIN_t(WX2615_t),
    .SDIN(CRC_OUT_8_28),
    .SDIN_t(CRC_OUT_8_28_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_29),
    .Q_t(CRC_OUT_8_29_t),
    .QN(n6096),
    .QN_t(n6096_t)
  );


  sdffs1
  \DFF_380/Q_reg 
  (
    .DIN(WX2613),
    .DIN_t(WX2613_t),
    .SDIN(CRC_OUT_8_27),
    .SDIN_t(CRC_OUT_8_27_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_28),
    .Q_t(CRC_OUT_8_28_t),
    .QN(n6087),
    .QN_t(n6087_t)
  );


  sdffs1
  \DFF_379/Q_reg 
  (
    .DIN(WX2611),
    .DIN_t(WX2611_t),
    .SDIN(CRC_OUT_8_26),
    .SDIN_t(CRC_OUT_8_26_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_27),
    .Q_t(CRC_OUT_8_27_t),
    .QN(n6078),
    .QN_t(n6078_t)
  );


  sdffs1
  \DFF_378/Q_reg 
  (
    .DIN(WX2609),
    .DIN_t(WX2609_t),
    .SDIN(CRC_OUT_8_25),
    .SDIN_t(CRC_OUT_8_25_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_26),
    .Q_t(CRC_OUT_8_26_t),
    .QN(n6069),
    .QN_t(n6069_t)
  );


  sdffs1
  \DFF_377/Q_reg 
  (
    .DIN(WX2607),
    .DIN_t(WX2607_t),
    .SDIN(CRC_OUT_8_24),
    .SDIN_t(CRC_OUT_8_24_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_25),
    .Q_t(CRC_OUT_8_25_t),
    .QN(n6060),
    .QN_t(n6060_t)
  );


  sdffs1
  \DFF_376/Q_reg 
  (
    .DIN(WX2605),
    .DIN_t(WX2605_t),
    .SDIN(CRC_OUT_8_23),
    .SDIN_t(CRC_OUT_8_23_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_24),
    .Q_t(CRC_OUT_8_24_t),
    .QN(n6051),
    .QN_t(n6051_t)
  );


  sdffs1
  \DFF_375/Q_reg 
  (
    .DIN(WX2603),
    .DIN_t(WX2603_t),
    .SDIN(CRC_OUT_8_22),
    .SDIN_t(CRC_OUT_8_22_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_23),
    .Q_t(CRC_OUT_8_23_t),
    .QN(n6042),
    .QN_t(n6042_t)
  );


  sdffs1
  \DFF_374/Q_reg 
  (
    .DIN(WX2601),
    .DIN_t(WX2601_t),
    .SDIN(CRC_OUT_8_21),
    .SDIN_t(CRC_OUT_8_21_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_22),
    .Q_t(CRC_OUT_8_22_t),
    .QN(n6033),
    .QN_t(n6033_t)
  );


  sdffs1
  \DFF_373/Q_reg 
  (
    .DIN(WX2599),
    .DIN_t(WX2599_t),
    .SDIN(CRC_OUT_8_20),
    .SDIN_t(CRC_OUT_8_20_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_21),
    .Q_t(CRC_OUT_8_21_t),
    .QN(n6024),
    .QN_t(n6024_t)
  );


  sdffs1
  \DFF_372/Q_reg 
  (
    .DIN(WX2597),
    .DIN_t(WX2597_t),
    .SDIN(CRC_OUT_8_19),
    .SDIN_t(CRC_OUT_8_19_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_20),
    .Q_t(CRC_OUT_8_20_t),
    .QN(n6015),
    .QN_t(n6015_t)
  );


  sdffs1
  \DFF_371/Q_reg 
  (
    .DIN(WX2595),
    .DIN_t(WX2595_t),
    .SDIN(CRC_OUT_8_18),
    .SDIN_t(CRC_OUT_8_18_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_19),
    .Q_t(CRC_OUT_8_19_t),
    .QN(n6006),
    .QN_t(n6006_t)
  );


  sdffs1
  \DFF_370/Q_reg 
  (
    .DIN(WX2593),
    .DIN_t(WX2593_t),
    .SDIN(CRC_OUT_8_17),
    .SDIN_t(CRC_OUT_8_17_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_18),
    .Q_t(CRC_OUT_8_18_t),
    .QN(n5997),
    .QN_t(n5997_t)
  );


  sdffs1
  \DFF_369/Q_reg 
  (
    .DIN(WX2591),
    .DIN_t(WX2591_t),
    .SDIN(CRC_OUT_8_16),
    .SDIN_t(CRC_OUT_8_16_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_17),
    .Q_t(CRC_OUT_8_17_t),
    .QN(n5988),
    .QN_t(n5988_t)
  );


  sdffs1
  \DFF_368/Q_reg 
  (
    .DIN(WX2589),
    .DIN_t(WX2589_t),
    .SDIN(CRC_OUT_8_15),
    .SDIN_t(CRC_OUT_8_15_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_16),
    .Q_t(CRC_OUT_8_16_t),
    .QN(n5979),
    .QN_t(n5979_t)
  );


  sdffs1
  \DFF_367/Q_reg 
  (
    .DIN(WX2587),
    .DIN_t(WX2587_t),
    .SDIN(CRC_OUT_8_14),
    .SDIN_t(CRC_OUT_8_14_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_15),
    .Q_t(CRC_OUT_8_15_t),
    .QN(n5970),
    .QN_t(n5970_t)
  );


  sdffs1
  \DFF_366/Q_reg 
  (
    .DIN(WX2585),
    .DIN_t(WX2585_t),
    .SDIN(CRC_OUT_8_13),
    .SDIN_t(CRC_OUT_8_13_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_14),
    .Q_t(CRC_OUT_8_14_t),
    .QN(n5963),
    .QN_t(n5963_t)
  );


  sdffs1
  \DFF_365/Q_reg 
  (
    .DIN(WX2583),
    .DIN_t(WX2583_t),
    .SDIN(CRC_OUT_8_12),
    .SDIN_t(CRC_OUT_8_12_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_13),
    .Q_t(CRC_OUT_8_13_t),
    .QN(n5956),
    .QN_t(n5956_t)
  );


  sdffs1
  \DFF_364/Q_reg 
  (
    .DIN(WX2581),
    .DIN_t(WX2581_t),
    .SDIN(CRC_OUT_8_11),
    .SDIN_t(CRC_OUT_8_11_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_12),
    .Q_t(CRC_OUT_8_12_t),
    .QN(n5949),
    .QN_t(n5949_t)
  );


  sdffs1
  \DFF_363/Q_reg 
  (
    .DIN(WX2579),
    .DIN_t(WX2579_t),
    .SDIN(CRC_OUT_8_10),
    .SDIN_t(CRC_OUT_8_10_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_11),
    .Q_t(CRC_OUT_8_11_t),
    .QN(n5942),
    .QN_t(n5942_t)
  );


  sdffs1
  \DFF_362/Q_reg 
  (
    .DIN(WX2577),
    .DIN_t(WX2577_t),
    .SDIN(CRC_OUT_8_9),
    .SDIN_t(CRC_OUT_8_9_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_10),
    .Q_t(CRC_OUT_8_10_t),
    .QN(n5935),
    .QN_t(n5935_t)
  );


  sdffs1
  \DFF_361/Q_reg 
  (
    .DIN(WX2575),
    .DIN_t(WX2575_t),
    .SDIN(CRC_OUT_8_8),
    .SDIN_t(CRC_OUT_8_8_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_9),
    .Q_t(CRC_OUT_8_9_t),
    .QN(n5928),
    .QN_t(n5928_t)
  );


  sdffs1
  \DFF_360/Q_reg 
  (
    .DIN(WX2573),
    .DIN_t(WX2573_t),
    .SDIN(CRC_OUT_8_7),
    .SDIN_t(CRC_OUT_8_7_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_8),
    .Q_t(CRC_OUT_8_8_t),
    .QN(n5921),
    .QN_t(n5921_t)
  );


  sdffs1
  \DFF_359/Q_reg 
  (
    .DIN(WX2571),
    .DIN_t(WX2571_t),
    .SDIN(CRC_OUT_8_6),
    .SDIN_t(CRC_OUT_8_6_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_7),
    .Q_t(CRC_OUT_8_7_t),
    .QN(n5914),
    .QN_t(n5914_t)
  );


  sdffs1
  \DFF_358/Q_reg 
  (
    .DIN(WX2569),
    .DIN_t(WX2569_t),
    .SDIN(CRC_OUT_8_5),
    .SDIN_t(CRC_OUT_8_5_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_6),
    .Q_t(CRC_OUT_8_6_t),
    .QN(n5907),
    .QN_t(n5907_t)
  );


  sdffs1
  \DFF_357/Q_reg 
  (
    .DIN(WX2567),
    .DIN_t(WX2567_t),
    .SDIN(CRC_OUT_8_4),
    .SDIN_t(CRC_OUT_8_4_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_5),
    .Q_t(CRC_OUT_8_5_t),
    .QN(n5900),
    .QN_t(n5900_t)
  );


  sdffs1
  \DFF_356/Q_reg 
  (
    .DIN(WX2565),
    .DIN_t(WX2565_t),
    .SDIN(CRC_OUT_8_3),
    .SDIN_t(CRC_OUT_8_3_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_4),
    .Q_t(CRC_OUT_8_4_t),
    .QN(n5893),
    .QN_t(n5893_t)
  );


  sdffs1
  \DFF_355/Q_reg 
  (
    .DIN(WX2563),
    .DIN_t(WX2563_t),
    .SDIN(CRC_OUT_8_2),
    .SDIN_t(CRC_OUT_8_2_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_3),
    .Q_t(CRC_OUT_8_3_t),
    .QN(n5886),
    .QN_t(n5886_t)
  );


  sdffs1
  \DFF_354/Q_reg 
  (
    .DIN(WX2561),
    .DIN_t(WX2561_t),
    .SDIN(CRC_OUT_8_1),
    .SDIN_t(CRC_OUT_8_1_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_2),
    .Q_t(CRC_OUT_8_2_t),
    .QN(n5879),
    .QN_t(n5879_t)
  );


  sdffs1
  \DFF_353/Q_reg 
  (
    .DIN(WX2559),
    .DIN_t(WX2559_t),
    .SDIN(CRC_OUT_8_0),
    .SDIN_t(CRC_OUT_8_0_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_1),
    .Q_t(CRC_OUT_8_1_t),
    .QN(n5872),
    .QN_t(n5872_t)
  );


  sdffs1
  \DFF_352/Q_reg 
  (
    .DIN(WX2557),
    .DIN_t(WX2557_t),
    .SDIN(n7098),
    .SDIN_t(n7098_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_8_0),
    .Q_t(CRC_OUT_8_0_t),
    .QN(n5865),
    .QN_t(n5865_t)
  );


  sdffs1
  \DFF_351/Q_reg 
  (
    .DIN(WX2191),
    .DIN_t(WX2191_t),
    .SDIN(n7097),
    .SDIN_t(n7097_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7098),
    .Q_t(n7098_t),
    .QN(n3286),
    .QN_t(n3286_t)
  );


  sdffs1
  \DFF_350/Q_reg 
  (
    .DIN(WX2189),
    .DIN_t(WX2189_t),
    .SDIN(n7096),
    .SDIN_t(n7096_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7097),
    .Q_t(n7097_t),
    .QN(n3288),
    .QN_t(n3288_t)
  );


  sdffs1
  \DFF_349/Q_reg 
  (
    .DIN(WX2187),
    .DIN_t(WX2187_t),
    .SDIN(n7095),
    .SDIN_t(n7095_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7096),
    .Q_t(n7096_t),
    .QN(n3290),
    .QN_t(n3290_t)
  );


  sdffs1
  \DFF_348/Q_reg 
  (
    .DIN(WX2185),
    .DIN_t(WX2185_t),
    .SDIN(n7094),
    .SDIN_t(n7094_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7095),
    .Q_t(n7095_t),
    .QN(n3292),
    .QN_t(n3292_t)
  );


  sdffs1
  \DFF_347/Q_reg 
  (
    .DIN(WX2183),
    .DIN_t(WX2183_t),
    .SDIN(n7093),
    .SDIN_t(n7093_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7094),
    .Q_t(n7094_t),
    .QN(n3294),
    .QN_t(n3294_t)
  );


  sdffs1
  \DFF_346/Q_reg 
  (
    .DIN(WX2181),
    .DIN_t(WX2181_t),
    .SDIN(n7092),
    .SDIN_t(n7092_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7093),
    .Q_t(n7093_t),
    .QN(n3296),
    .QN_t(n3296_t)
  );


  sdffs1
  \DFF_345/Q_reg 
  (
    .DIN(WX2179),
    .DIN_t(WX2179_t),
    .SDIN(n7091),
    .SDIN_t(n7091_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7092),
    .Q_t(n7092_t),
    .QN(n3298),
    .QN_t(n3298_t)
  );


  sdffs1
  \DFF_344/Q_reg 
  (
    .DIN(WX2177),
    .DIN_t(WX2177_t),
    .SDIN(n7090),
    .SDIN_t(n7090_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7091),
    .Q_t(n7091_t),
    .QN(n3300),
    .QN_t(n3300_t)
  );


  sdffs1
  \DFF_343/Q_reg 
  (
    .DIN(WX2175),
    .DIN_t(WX2175_t),
    .SDIN(n7089),
    .SDIN_t(n7089_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7090),
    .Q_t(n7090_t),
    .QN(n3302),
    .QN_t(n3302_t)
  );


  sdffs1
  \DFF_342/Q_reg 
  (
    .DIN(WX2173),
    .DIN_t(WX2173_t),
    .SDIN(n7088),
    .SDIN_t(n7088_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7089),
    .Q_t(n7089_t),
    .QN(n3304),
    .QN_t(n3304_t)
  );


  sdffs1
  \DFF_341/Q_reg 
  (
    .DIN(WX2171),
    .DIN_t(WX2171_t),
    .SDIN(n7087),
    .SDIN_t(n7087_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7088),
    .Q_t(n7088_t),
    .QN(n3306),
    .QN_t(n3306_t)
  );


  sdffs1
  \DFF_340/Q_reg 
  (
    .DIN(WX2169),
    .DIN_t(WX2169_t),
    .SDIN(n7086),
    .SDIN_t(n7086_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7087),
    .Q_t(n7087_t),
    .QN(n3308),
    .QN_t(n3308_t)
  );


  sdffs1
  \DFF_339/Q_reg 
  (
    .DIN(WX2167),
    .DIN_t(WX2167_t),
    .SDIN(n7085),
    .SDIN_t(n7085_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7086),
    .Q_t(n7086_t),
    .QN(n3310),
    .QN_t(n3310_t)
  );


  sdffs1
  \DFF_338/Q_reg 
  (
    .DIN(WX2165),
    .DIN_t(WX2165_t),
    .SDIN(n7084),
    .SDIN_t(n7084_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7085),
    .Q_t(n7085_t),
    .QN(n3312),
    .QN_t(n3312_t)
  );


  sdffs1
  \DFF_337/Q_reg 
  (
    .DIN(WX2163),
    .DIN_t(WX2163_t),
    .SDIN(n7083),
    .SDIN_t(n7083_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7084),
    .Q_t(n7084_t),
    .QN(n3314),
    .QN_t(n3314_t)
  );


  sdffs1
  \DFF_336/Q_reg 
  (
    .DIN(WX2161),
    .DIN_t(WX2161_t),
    .SDIN(n7082),
    .SDIN_t(n7082_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7083),
    .Q_t(n7083_t),
    .QN(n3316),
    .QN_t(n3316_t)
  );


  sdffs1
  \DFF_335/Q_reg 
  (
    .DIN(WX2159),
    .DIN_t(WX2159_t),
    .SDIN(n7081),
    .SDIN_t(n7081_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7082),
    .Q_t(n7082_t),
    .QN(n5978),
    .QN_t(n5978_t)
  );


  sdffs1
  \DFF_334/Q_reg 
  (
    .DIN(WX2157),
    .DIN_t(WX2157_t),
    .SDIN(n7080),
    .SDIN_t(n7080_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7081),
    .Q_t(n7081_t),
    .QN(n5987),
    .QN_t(n5987_t)
  );


  sdffs1
  \DFF_333/Q_reg 
  (
    .DIN(WX2155),
    .DIN_t(WX2155_t),
    .SDIN(n7079),
    .SDIN_t(n7079_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7080),
    .Q_t(n7080_t),
    .QN(n5996),
    .QN_t(n5996_t)
  );


  sdffs1
  \DFF_332/Q_reg 
  (
    .DIN(WX2153),
    .DIN_t(WX2153_t),
    .SDIN(n7078),
    .SDIN_t(n7078_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7079),
    .Q_t(n7079_t),
    .QN(n6005),
    .QN_t(n6005_t)
  );


  sdffs1
  \DFF_331/Q_reg 
  (
    .DIN(WX2151),
    .DIN_t(WX2151_t),
    .SDIN(n7077),
    .SDIN_t(n7077_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7078),
    .Q_t(n7078_t),
    .QN(n6014),
    .QN_t(n6014_t)
  );


  sdffs1
  \DFF_330/Q_reg 
  (
    .DIN(WX2149),
    .DIN_t(WX2149_t),
    .SDIN(n7076),
    .SDIN_t(n7076_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7077),
    .Q_t(n7077_t),
    .QN(n6023),
    .QN_t(n6023_t)
  );


  sdffs1
  \DFF_329/Q_reg 
  (
    .DIN(WX2147),
    .DIN_t(WX2147_t),
    .SDIN(n7075),
    .SDIN_t(n7075_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7076),
    .Q_t(n7076_t),
    .QN(n6032),
    .QN_t(n6032_t)
  );


  sdffs1
  \DFF_328/Q_reg 
  (
    .DIN(WX2145),
    .DIN_t(WX2145_t),
    .SDIN(n7074),
    .SDIN_t(n7074_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7075),
    .Q_t(n7075_t),
    .QN(n6041),
    .QN_t(n6041_t)
  );


  sdffs1
  \DFF_327/Q_reg 
  (
    .DIN(WX2143),
    .DIN_t(WX2143_t),
    .SDIN(n7073),
    .SDIN_t(n7073_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7074),
    .Q_t(n7074_t),
    .QN(n6050),
    .QN_t(n6050_t)
  );


  sdffs1
  \DFF_326/Q_reg 
  (
    .DIN(WX2141),
    .DIN_t(WX2141_t),
    .SDIN(n7072),
    .SDIN_t(n7072_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7073),
    .Q_t(n7073_t),
    .QN(n6059),
    .QN_t(n6059_t)
  );


  sdffs1
  \DFF_325/Q_reg 
  (
    .DIN(WX2139),
    .DIN_t(WX2139_t),
    .SDIN(n7071),
    .SDIN_t(n7071_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7072),
    .Q_t(n7072_t),
    .QN(n6068),
    .QN_t(n6068_t)
  );


  sdffs1
  \DFF_324/Q_reg 
  (
    .DIN(WX2137),
    .DIN_t(WX2137_t),
    .SDIN(n7070),
    .SDIN_t(n7070_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7071),
    .Q_t(n7071_t),
    .QN(n6077),
    .QN_t(n6077_t)
  );


  sdffs1
  \DFF_323/Q_reg 
  (
    .DIN(WX2135),
    .DIN_t(WX2135_t),
    .SDIN(n7069),
    .SDIN_t(n7069_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7070),
    .Q_t(n7070_t),
    .QN(n6086),
    .QN_t(n6086_t)
  );


  sdffs1
  \DFF_322/Q_reg 
  (
    .DIN(WX2133),
    .DIN_t(WX2133_t),
    .SDIN(n7068),
    .SDIN_t(n7068_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7069),
    .Q_t(n7069_t),
    .QN(n6095),
    .QN_t(n6095_t)
  );


  sdffs1
  \DFF_321/Q_reg 
  (
    .DIN(WX2131),
    .DIN_t(WX2131_t),
    .SDIN(n7067),
    .SDIN_t(n7067_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7068),
    .Q_t(n7068_t),
    .QN(n6104),
    .QN_t(n6104_t)
  );


  sdffs1
  \DFF_320/Q_reg 
  (
    .DIN(WX2129),
    .DIN_t(WX2129_t),
    .SDIN(n7066),
    .SDIN_t(n7066_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7067),
    .Q_t(n7067_t),
    .QN(n6113),
    .QN_t(n6113_t)
  );


  sdffs1
  \DFF_319/Q_reg 
  (
    .DIN(WX2127),
    .DIN_t(WX2127_t),
    .SDIN(n7065),
    .SDIN_t(n7065_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7066),
    .Q_t(n7066_t),
    .QN(n5864),
    .QN_t(n5864_t)
  );


  sdffs1
  \DFF_318/Q_reg 
  (
    .DIN(WX2125),
    .DIN_t(WX2125_t),
    .SDIN(n7064),
    .SDIN_t(n7064_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7065),
    .Q_t(n7065_t),
    .QN(n5871),
    .QN_t(n5871_t)
  );


  sdffs1
  \DFF_317/Q_reg 
  (
    .DIN(WX2123),
    .DIN_t(WX2123_t),
    .SDIN(n7063),
    .SDIN_t(n7063_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7064),
    .Q_t(n7064_t),
    .QN(n5878),
    .QN_t(n5878_t)
  );


  sdffs1
  \DFF_316/Q_reg 
  (
    .DIN(WX2121),
    .DIN_t(WX2121_t),
    .SDIN(n7062),
    .SDIN_t(n7062_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7063),
    .Q_t(n7063_t),
    .QN(n5885),
    .QN_t(n5885_t)
  );


  sdffs1
  \DFF_315/Q_reg 
  (
    .DIN(WX2119),
    .DIN_t(WX2119_t),
    .SDIN(n7061),
    .SDIN_t(n7061_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7062),
    .Q_t(n7062_t),
    .QN(n5892),
    .QN_t(n5892_t)
  );


  sdffs1
  \DFF_314/Q_reg 
  (
    .DIN(WX2117),
    .DIN_t(WX2117_t),
    .SDIN(n7060),
    .SDIN_t(n7060_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7061),
    .Q_t(n7061_t),
    .QN(n5899),
    .QN_t(n5899_t)
  );


  sdffs1
  \DFF_313/Q_reg 
  (
    .DIN(WX2115),
    .DIN_t(WX2115_t),
    .SDIN(n7059),
    .SDIN_t(n7059_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7060),
    .Q_t(n7060_t),
    .QN(n5906),
    .QN_t(n5906_t)
  );


  sdffs1
  \DFF_312/Q_reg 
  (
    .DIN(WX2113),
    .DIN_t(WX2113_t),
    .SDIN(n7058),
    .SDIN_t(n7058_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7059),
    .Q_t(n7059_t),
    .QN(n5913),
    .QN_t(n5913_t)
  );


  sdffs1
  \DFF_311/Q_reg 
  (
    .DIN(WX2111),
    .DIN_t(WX2111_t),
    .SDIN(n7057),
    .SDIN_t(n7057_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7058),
    .Q_t(n7058_t),
    .QN(n5920),
    .QN_t(n5920_t)
  );


  sdffs1
  \DFF_310/Q_reg 
  (
    .DIN(WX2109),
    .DIN_t(WX2109_t),
    .SDIN(n7056),
    .SDIN_t(n7056_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7057),
    .Q_t(n7057_t),
    .QN(n5927),
    .QN_t(n5927_t)
  );


  sdffs1
  \DFF_309/Q_reg 
  (
    .DIN(WX2107),
    .DIN_t(WX2107_t),
    .SDIN(n7055),
    .SDIN_t(n7055_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7056),
    .Q_t(n7056_t),
    .QN(n5934),
    .QN_t(n5934_t)
  );


  sdffs1
  \DFF_308/Q_reg 
  (
    .DIN(WX2105),
    .DIN_t(WX2105_t),
    .SDIN(n7054),
    .SDIN_t(n7054_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7055),
    .Q_t(n7055_t),
    .QN(n5941),
    .QN_t(n5941_t)
  );


  sdffs1
  \DFF_307/Q_reg 
  (
    .DIN(WX2103),
    .DIN_t(WX2103_t),
    .SDIN(n7053),
    .SDIN_t(n7053_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7054),
    .Q_t(n7054_t),
    .QN(n5948),
    .QN_t(n5948_t)
  );


  sdffs1
  \DFF_306/Q_reg 
  (
    .DIN(WX2101),
    .DIN_t(WX2101_t),
    .SDIN(n7052),
    .SDIN_t(n7052_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7053),
    .Q_t(n7053_t),
    .QN(n5955),
    .QN_t(n5955_t)
  );


  sdffs1
  \DFF_305/Q_reg 
  (
    .DIN(WX2099),
    .DIN_t(WX2099_t),
    .SDIN(n7051),
    .SDIN_t(n7051_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7052),
    .Q_t(n7052_t),
    .QN(n5962),
    .QN_t(n5962_t)
  );


  sdffs1
  \DFF_304/Q_reg 
  (
    .DIN(WX2097),
    .DIN_t(WX2097_t),
    .SDIN(n7050),
    .SDIN_t(n7050_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7051),
    .Q_t(n7051_t),
    .QN(n5969),
    .QN_t(n5969_t)
  );


  sdffs1
  \DFF_303/Q_reg 
  (
    .DIN(WX2095),
    .DIN_t(WX2095_t),
    .SDIN(n7049),
    .SDIN_t(n7049_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7050),
    .Q_t(n7050_t),
    .QN(n5977),
    .QN_t(n5977_t)
  );


  sdffs1
  \DFF_302/Q_reg 
  (
    .DIN(WX2093),
    .DIN_t(WX2093_t),
    .SDIN(n7048),
    .SDIN_t(n7048_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7049),
    .Q_t(n7049_t),
    .QN(n5986),
    .QN_t(n5986_t)
  );


  sdffs1
  \DFF_301/Q_reg 
  (
    .DIN(WX2091),
    .DIN_t(WX2091_t),
    .SDIN(n7047),
    .SDIN_t(n7047_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7048),
    .Q_t(n7048_t),
    .QN(n5995),
    .QN_t(n5995_t)
  );


  sdffs1
  \DFF_300/Q_reg 
  (
    .DIN(WX2089),
    .DIN_t(WX2089_t),
    .SDIN(n7046),
    .SDIN_t(n7046_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7047),
    .Q_t(n7047_t),
    .QN(n6004),
    .QN_t(n6004_t)
  );


  sdffs1
  \DFF_299/Q_reg 
  (
    .DIN(WX2087),
    .DIN_t(WX2087_t),
    .SDIN(n7045),
    .SDIN_t(n7045_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7046),
    .Q_t(n7046_t),
    .QN(n6013),
    .QN_t(n6013_t)
  );


  sdffs1
  \DFF_298/Q_reg 
  (
    .DIN(WX2085),
    .DIN_t(WX2085_t),
    .SDIN(n7044),
    .SDIN_t(n7044_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7045),
    .Q_t(n7045_t),
    .QN(n6022),
    .QN_t(n6022_t)
  );


  sdffs1
  \DFF_297/Q_reg 
  (
    .DIN(WX2083),
    .DIN_t(WX2083_t),
    .SDIN(n7043),
    .SDIN_t(n7043_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7044),
    .Q_t(n7044_t),
    .QN(n6031),
    .QN_t(n6031_t)
  );


  sdffs1
  \DFF_296/Q_reg 
  (
    .DIN(WX2081),
    .DIN_t(WX2081_t),
    .SDIN(n7042),
    .SDIN_t(n7042_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7043),
    .Q_t(n7043_t),
    .QN(n6040),
    .QN_t(n6040_t)
  );


  sdffs1
  \DFF_295/Q_reg 
  (
    .DIN(WX2079),
    .DIN_t(WX2079_t),
    .SDIN(n7041),
    .SDIN_t(n7041_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7042),
    .Q_t(n7042_t),
    .QN(n6049),
    .QN_t(n6049_t)
  );


  sdffs1
  \DFF_294/Q_reg 
  (
    .DIN(WX2077),
    .DIN_t(WX2077_t),
    .SDIN(n7040),
    .SDIN_t(n7040_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7041),
    .Q_t(n7041_t),
    .QN(n6058),
    .QN_t(n6058_t)
  );


  sdffs1
  \DFF_293/Q_reg 
  (
    .DIN(WX2075),
    .DIN_t(WX2075_t),
    .SDIN(n7039),
    .SDIN_t(n7039_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7040),
    .Q_t(n7040_t),
    .QN(n6067),
    .QN_t(n6067_t)
  );


  sdffs1
  \DFF_292/Q_reg 
  (
    .DIN(WX2073),
    .DIN_t(WX2073_t),
    .SDIN(n7038),
    .SDIN_t(n7038_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7039),
    .Q_t(n7039_t),
    .QN(n6076),
    .QN_t(n6076_t)
  );


  sdffs1
  \DFF_291/Q_reg 
  (
    .DIN(WX2071),
    .DIN_t(WX2071_t),
    .SDIN(n7037),
    .SDIN_t(n7037_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7038),
    .Q_t(n7038_t),
    .QN(n6085),
    .QN_t(n6085_t)
  );


  sdffs1
  \DFF_290/Q_reg 
  (
    .DIN(WX2069),
    .DIN_t(WX2069_t),
    .SDIN(n7036),
    .SDIN_t(n7036_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7037),
    .Q_t(n7037_t),
    .QN(n6094),
    .QN_t(n6094_t)
  );


  sdffs1
  \DFF_289/Q_reg 
  (
    .DIN(WX2067),
    .DIN_t(WX2067_t),
    .SDIN(n7035),
    .SDIN_t(n7035_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7036),
    .Q_t(n7036_t),
    .QN(n6103),
    .QN_t(n6103_t)
  );


  sdffs1
  \DFF_288/Q_reg 
  (
    .DIN(WX2065),
    .DIN_t(WX2065_t),
    .SDIN(n5863),
    .SDIN_t(n5863_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7035),
    .Q_t(n7035_t),
    .QN(n6112),
    .QN_t(n6112_t)
  );


  sdffs1
  \DFF_287/Q_reg 
  (
    .DIN(WX2063),
    .DIN_t(WX2063_t),
    .SDIN(n5870),
    .SDIN_t(n5870_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5863),
    .Q_t(n5863_t)
  );


  sdffs1
  \DFF_286/Q_reg 
  (
    .DIN(WX2061),
    .DIN_t(WX2061_t),
    .SDIN(n5877),
    .SDIN_t(n5877_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5870),
    .Q_t(n5870_t)
  );


  sdffs1
  \DFF_285/Q_reg 
  (
    .DIN(WX2059),
    .DIN_t(WX2059_t),
    .SDIN(n5884),
    .SDIN_t(n5884_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5877),
    .Q_t(n5877_t)
  );


  sdffs1
  \DFF_284/Q_reg 
  (
    .DIN(WX2057),
    .DIN_t(WX2057_t),
    .SDIN(n5891),
    .SDIN_t(n5891_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5884),
    .Q_t(n5884_t)
  );


  sdffs1
  \DFF_283/Q_reg 
  (
    .DIN(WX2055),
    .DIN_t(WX2055_t),
    .SDIN(n5898),
    .SDIN_t(n5898_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5891),
    .Q_t(n5891_t)
  );


  sdffs1
  \DFF_282/Q_reg 
  (
    .DIN(WX2053),
    .DIN_t(WX2053_t),
    .SDIN(n5905),
    .SDIN_t(n5905_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5898),
    .Q_t(n5898_t)
  );


  sdffs1
  \DFF_281/Q_reg 
  (
    .DIN(WX2051),
    .DIN_t(WX2051_t),
    .SDIN(n5912),
    .SDIN_t(n5912_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5905),
    .Q_t(n5905_t)
  );


  sdffs1
  \DFF_280/Q_reg 
  (
    .DIN(WX2049),
    .DIN_t(WX2049_t),
    .SDIN(n5919),
    .SDIN_t(n5919_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5912),
    .Q_t(n5912_t)
  );


  sdffs1
  \DFF_279/Q_reg 
  (
    .DIN(WX2047),
    .DIN_t(WX2047_t),
    .SDIN(n5926),
    .SDIN_t(n5926_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5919),
    .Q_t(n5919_t)
  );


  sdffs1
  \DFF_278/Q_reg 
  (
    .DIN(WX2045),
    .DIN_t(WX2045_t),
    .SDIN(n5933),
    .SDIN_t(n5933_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5926),
    .Q_t(n5926_t)
  );


  sdffs1
  \DFF_277/Q_reg 
  (
    .DIN(WX2043),
    .DIN_t(WX2043_t),
    .SDIN(n5940),
    .SDIN_t(n5940_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5933),
    .Q_t(n5933_t)
  );


  sdffs1
  \DFF_276/Q_reg 
  (
    .DIN(WX2041),
    .DIN_t(WX2041_t),
    .SDIN(n5947),
    .SDIN_t(n5947_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5940),
    .Q_t(n5940_t)
  );


  sdffs1
  \DFF_275/Q_reg 
  (
    .DIN(WX2039),
    .DIN_t(WX2039_t),
    .SDIN(n5954),
    .SDIN_t(n5954_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5947),
    .Q_t(n5947_t)
  );


  sdffs1
  \DFF_274/Q_reg 
  (
    .DIN(WX2037),
    .DIN_t(WX2037_t),
    .SDIN(n5961),
    .SDIN_t(n5961_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5954),
    .Q_t(n5954_t)
  );


  sdffs1
  \DFF_273/Q_reg 
  (
    .DIN(WX2035),
    .DIN_t(WX2035_t),
    .SDIN(n5968),
    .SDIN_t(n5968_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5961),
    .Q_t(n5961_t)
  );


  sdffs1
  \DFF_272/Q_reg 
  (
    .DIN(WX2033),
    .DIN_t(WX2033_t),
    .SDIN(n5976),
    .SDIN_t(n5976_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5968),
    .Q_t(n5968_t)
  );


  sdffs1
  \DFF_271/Q_reg 
  (
    .DIN(WX2031),
    .DIN_t(WX2031_t),
    .SDIN(n5985),
    .SDIN_t(n5985_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5976),
    .Q_t(n5976_t)
  );


  sdffs1
  \DFF_270/Q_reg 
  (
    .DIN(WX2029),
    .DIN_t(WX2029_t),
    .SDIN(n5994),
    .SDIN_t(n5994_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5985),
    .Q_t(n5985_t)
  );


  sdffs1
  \DFF_269/Q_reg 
  (
    .DIN(WX2027),
    .DIN_t(WX2027_t),
    .SDIN(n6003),
    .SDIN_t(n6003_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n5994),
    .Q_t(n5994_t)
  );


  sdffs1
  \DFF_268/Q_reg 
  (
    .DIN(WX2025),
    .DIN_t(WX2025_t),
    .SDIN(n6012),
    .SDIN_t(n6012_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6003),
    .Q_t(n6003_t)
  );


  sdffs1
  \DFF_267/Q_reg 
  (
    .DIN(WX2023),
    .DIN_t(WX2023_t),
    .SDIN(n6021),
    .SDIN_t(n6021_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6012),
    .Q_t(n6012_t)
  );


  sdffs1
  \DFF_266/Q_reg 
  (
    .DIN(WX2021),
    .DIN_t(WX2021_t),
    .SDIN(n6030),
    .SDIN_t(n6030_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6021),
    .Q_t(n6021_t)
  );


  sdffs1
  \DFF_265/Q_reg 
  (
    .DIN(WX2019),
    .DIN_t(WX2019_t),
    .SDIN(n6039),
    .SDIN_t(n6039_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6030),
    .Q_t(n6030_t)
  );


  sdffs1
  \DFF_264/Q_reg 
  (
    .DIN(WX2017),
    .DIN_t(WX2017_t),
    .SDIN(n6048),
    .SDIN_t(n6048_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6039),
    .Q_t(n6039_t)
  );


  sdffs1
  \DFF_263/Q_reg 
  (
    .DIN(WX2015),
    .DIN_t(WX2015_t),
    .SDIN(n6057),
    .SDIN_t(n6057_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6048),
    .Q_t(n6048_t)
  );


  sdffs1
  \DFF_262/Q_reg 
  (
    .DIN(WX2013),
    .DIN_t(WX2013_t),
    .SDIN(n6066),
    .SDIN_t(n6066_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6057),
    .Q_t(n6057_t)
  );


  sdffs1
  \DFF_261/Q_reg 
  (
    .DIN(WX2011),
    .DIN_t(WX2011_t),
    .SDIN(n6075),
    .SDIN_t(n6075_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6066),
    .Q_t(n6066_t)
  );


  sdffs1
  \DFF_260/Q_reg 
  (
    .DIN(WX2009),
    .DIN_t(WX2009_t),
    .SDIN(n6084),
    .SDIN_t(n6084_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6075),
    .Q_t(n6075_t)
  );


  sdffs1
  \DFF_259/Q_reg 
  (
    .DIN(WX2007),
    .DIN_t(WX2007_t),
    .SDIN(n6093),
    .SDIN_t(n6093_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6084),
    .Q_t(n6084_t)
  );


  sdffs1
  \DFF_258/Q_reg 
  (
    .DIN(WX2005),
    .DIN_t(WX2005_t),
    .SDIN(n6102),
    .SDIN_t(n6102_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6093),
    .Q_t(n6093_t)
  );


  sdffs1
  \DFF_257/Q_reg 
  (
    .DIN(WX2003),
    .DIN_t(WX2003_t),
    .SDIN(n6111),
    .SDIN_t(n6111_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6102),
    .Q_t(n6102_t)
  );


  sdffs1
  \DFF_256/Q_reg 
  (
    .DIN(WX2001),
    .DIN_t(WX2001_t),
    .SDIN(n7034),
    .SDIN_t(n7034_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6111),
    .Q_t(n6111_t)
  );


  sdffs1
  \DFF_255/Q_reg 
  (
    .DIN(WX1999),
    .DIN_t(WX1999_t),
    .SDIN(n7033),
    .SDIN_t(n7033_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7034),
    .Q_t(n7034_t),
    .QN(n5862),
    .QN_t(n5862_t)
  );


  sdffs1
  \DFF_254/Q_reg 
  (
    .DIN(WX1997),
    .DIN_t(WX1997_t),
    .SDIN(n7032),
    .SDIN_t(n7032_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7033),
    .Q_t(n7033_t),
    .QN(n5869),
    .QN_t(n5869_t)
  );


  sdffs1
  \DFF_253/Q_reg 
  (
    .DIN(WX1995),
    .DIN_t(WX1995_t),
    .SDIN(n7031),
    .SDIN_t(n7031_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7032),
    .Q_t(n7032_t),
    .QN(n5876),
    .QN_t(n5876_t)
  );


  sdffs1
  \DFF_252/Q_reg 
  (
    .DIN(WX1993),
    .DIN_t(WX1993_t),
    .SDIN(n7030),
    .SDIN_t(n7030_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7031),
    .Q_t(n7031_t),
    .QN(n5883),
    .QN_t(n5883_t)
  );


  sdffs1
  \DFF_251/Q_reg 
  (
    .DIN(WX1991),
    .DIN_t(WX1991_t),
    .SDIN(n7029),
    .SDIN_t(n7029_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7030),
    .Q_t(n7030_t),
    .QN(n5890),
    .QN_t(n5890_t)
  );


  sdffs1
  \DFF_250/Q_reg 
  (
    .DIN(WX1989),
    .DIN_t(WX1989_t),
    .SDIN(n7028),
    .SDIN_t(n7028_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7029),
    .Q_t(n7029_t),
    .QN(n5897),
    .QN_t(n5897_t)
  );


  sdffs1
  \DFF_249/Q_reg 
  (
    .DIN(WX1987),
    .DIN_t(WX1987_t),
    .SDIN(n7027),
    .SDIN_t(n7027_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7028),
    .Q_t(n7028_t),
    .QN(n5904),
    .QN_t(n5904_t)
  );


  sdffs1
  \DFF_248/Q_reg 
  (
    .DIN(WX1985),
    .DIN_t(WX1985_t),
    .SDIN(n7026),
    .SDIN_t(n7026_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7027),
    .Q_t(n7027_t),
    .QN(n5911),
    .QN_t(n5911_t)
  );


  sdffs1
  \DFF_247/Q_reg 
  (
    .DIN(WX1983),
    .DIN_t(WX1983_t),
    .SDIN(n7025),
    .SDIN_t(n7025_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7026),
    .Q_t(n7026_t),
    .QN(n5918),
    .QN_t(n5918_t)
  );


  sdffs1
  \DFF_246/Q_reg 
  (
    .DIN(WX1981),
    .DIN_t(WX1981_t),
    .SDIN(n7024),
    .SDIN_t(n7024_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7025),
    .Q_t(n7025_t),
    .QN(n5925),
    .QN_t(n5925_t)
  );


  sdffs1
  \DFF_245/Q_reg 
  (
    .DIN(WX1979),
    .DIN_t(WX1979_t),
    .SDIN(n7023),
    .SDIN_t(n7023_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7024),
    .Q_t(n7024_t),
    .QN(n5932),
    .QN_t(n5932_t)
  );


  sdffs1
  \DFF_244/Q_reg 
  (
    .DIN(WX1977),
    .DIN_t(WX1977_t),
    .SDIN(n7022),
    .SDIN_t(n7022_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7023),
    .Q_t(n7023_t),
    .QN(n5939),
    .QN_t(n5939_t)
  );


  sdffs1
  \DFF_243/Q_reg 
  (
    .DIN(WX1975),
    .DIN_t(WX1975_t),
    .SDIN(n7021),
    .SDIN_t(n7021_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7022),
    .Q_t(n7022_t),
    .QN(n5946),
    .QN_t(n5946_t)
  );


  sdffs1
  \DFF_242/Q_reg 
  (
    .DIN(WX1973),
    .DIN_t(WX1973_t),
    .SDIN(n7020),
    .SDIN_t(n7020_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7021),
    .Q_t(n7021_t),
    .QN(n5953),
    .QN_t(n5953_t)
  );


  sdffs1
  \DFF_241/Q_reg 
  (
    .DIN(WX1971),
    .DIN_t(WX1971_t),
    .SDIN(n7019),
    .SDIN_t(n7019_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7020),
    .Q_t(n7020_t),
    .QN(n5960),
    .QN_t(n5960_t)
  );


  sdffs1
  \DFF_240/Q_reg 
  (
    .DIN(WX1969),
    .DIN_t(WX1969_t),
    .SDIN(n7018),
    .SDIN_t(n7018_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7019),
    .Q_t(n7019_t),
    .QN(n5967),
    .QN_t(n5967_t)
  );


  sdffs1
  \DFF_239/Q_reg 
  (
    .DIN(WX1967),
    .DIN_t(WX1967_t),
    .SDIN(n7017),
    .SDIN_t(n7017_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7018),
    .Q_t(n7018_t),
    .QN(n5975),
    .QN_t(n5975_t)
  );


  sdffs1
  \DFF_238/Q_reg 
  (
    .DIN(WX1965),
    .DIN_t(WX1965_t),
    .SDIN(n7016),
    .SDIN_t(n7016_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7017),
    .Q_t(n7017_t),
    .QN(n5984),
    .QN_t(n5984_t)
  );


  sdffs1
  \DFF_237/Q_reg 
  (
    .DIN(WX1963),
    .DIN_t(WX1963_t),
    .SDIN(n7015),
    .SDIN_t(n7015_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7016),
    .Q_t(n7016_t),
    .QN(n5993),
    .QN_t(n5993_t)
  );


  sdffs1
  \DFF_236/Q_reg 
  (
    .DIN(WX1961),
    .DIN_t(WX1961_t),
    .SDIN(n7014),
    .SDIN_t(n7014_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7015),
    .Q_t(n7015_t),
    .QN(n6002),
    .QN_t(n6002_t)
  );


  sdffs1
  \DFF_235/Q_reg 
  (
    .DIN(WX1959),
    .DIN_t(WX1959_t),
    .SDIN(n7013),
    .SDIN_t(n7013_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7014),
    .Q_t(n7014_t),
    .QN(n6011),
    .QN_t(n6011_t)
  );


  sdffs1
  \DFF_234/Q_reg 
  (
    .DIN(WX1957),
    .DIN_t(WX1957_t),
    .SDIN(n7012),
    .SDIN_t(n7012_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7013),
    .Q_t(n7013_t),
    .QN(n6020),
    .QN_t(n6020_t)
  );


  sdffs1
  \DFF_233/Q_reg 
  (
    .DIN(WX1955),
    .DIN_t(WX1955_t),
    .SDIN(n7011),
    .SDIN_t(n7011_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7012),
    .Q_t(n7012_t),
    .QN(n6029),
    .QN_t(n6029_t)
  );


  sdffs1
  \DFF_232/Q_reg 
  (
    .DIN(WX1953),
    .DIN_t(WX1953_t),
    .SDIN(n7010),
    .SDIN_t(n7010_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7011),
    .Q_t(n7011_t),
    .QN(n6038),
    .QN_t(n6038_t)
  );


  sdffs1
  \DFF_231/Q_reg 
  (
    .DIN(WX1951),
    .DIN_t(WX1951_t),
    .SDIN(n7009),
    .SDIN_t(n7009_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7010),
    .Q_t(n7010_t),
    .QN(n6047),
    .QN_t(n6047_t)
  );


  sdffs1
  \DFF_230/Q_reg 
  (
    .DIN(WX1949),
    .DIN_t(WX1949_t),
    .SDIN(n7008),
    .SDIN_t(n7008_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7009),
    .Q_t(n7009_t),
    .QN(n6056),
    .QN_t(n6056_t)
  );


  sdffs1
  \DFF_229/Q_reg 
  (
    .DIN(WX1947),
    .DIN_t(WX1947_t),
    .SDIN(n7007),
    .SDIN_t(n7007_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7008),
    .Q_t(n7008_t),
    .QN(n6065),
    .QN_t(n6065_t)
  );


  sdffs1
  \DFF_228/Q_reg 
  (
    .DIN(WX1945),
    .DIN_t(WX1945_t),
    .SDIN(n7006),
    .SDIN_t(n7006_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7007),
    .Q_t(n7007_t),
    .QN(n6074),
    .QN_t(n6074_t)
  );


  sdffs1
  \DFF_227/Q_reg 
  (
    .DIN(WX1943),
    .DIN_t(WX1943_t),
    .SDIN(n7005),
    .SDIN_t(n7005_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7006),
    .Q_t(n7006_t),
    .QN(n6083),
    .QN_t(n6083_t)
  );


  sdffs1
  \DFF_226/Q_reg 
  (
    .DIN(WX1941),
    .DIN_t(WX1941_t),
    .SDIN(n7004),
    .SDIN_t(n7004_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7005),
    .Q_t(n7005_t),
    .QN(n6092),
    .QN_t(n6092_t)
  );


  sdffs1
  \DFF_225/Q_reg 
  (
    .DIN(WX1939),
    .DIN_t(WX1939_t),
    .SDIN(n7003),
    .SDIN_t(n7003_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7004),
    .Q_t(n7004_t),
    .QN(n6101),
    .QN_t(n6101_t)
  );


  sdffs1
  \DFF_224/Q_reg 
  (
    .DIN(WX1937),
    .DIN_t(WX1937_t),
    .SDIN(n7002),
    .SDIN_t(n7002_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7003),
    .Q_t(n7003_t),
    .QN(n6110),
    .QN_t(n6110_t)
  );


  sdffs1
  \DFF_223/Q_reg 
  (
    .DIN(WX1839),
    .DIN_t(WX1839_t),
    .SDIN(n7001),
    .SDIN_t(n7001_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7002),
    .Q_t(n7002_t),
    .QN(n6116),
    .QN_t(n6116_t)
  );


  sdffs1
  \DFF_222/Q_reg 
  (
    .DIN(WX1837),
    .DIN_t(WX1837_t),
    .SDIN(n7000),
    .SDIN_t(n7000_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7001),
    .Q_t(n7001_t),
    .QN(n6117),
    .QN_t(n6117_t)
  );


  sdffs1
  \DFF_221/Q_reg 
  (
    .DIN(WX1835),
    .DIN_t(WX1835_t),
    .SDIN(n6999),
    .SDIN_t(n6999_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n7000),
    .Q_t(n7000_t),
    .QN(n6118),
    .QN_t(n6118_t)
  );


  sdffs1
  \DFF_220/Q_reg 
  (
    .DIN(WX1833),
    .DIN_t(WX1833_t),
    .SDIN(n6998),
    .SDIN_t(n6998_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6999),
    .Q_t(n6999_t),
    .QN(n6119),
    .QN_t(n6119_t)
  );


  sdffs1
  \DFF_219/Q_reg 
  (
    .DIN(WX1831),
    .DIN_t(WX1831_t),
    .SDIN(n6997),
    .SDIN_t(n6997_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6998),
    .Q_t(n6998_t),
    .QN(n6120),
    .QN_t(n6120_t)
  );


  sdffs1
  \DFF_218/Q_reg 
  (
    .DIN(WX1829),
    .DIN_t(WX1829_t),
    .SDIN(n6996),
    .SDIN_t(n6996_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6997),
    .Q_t(n6997_t),
    .QN(n6121),
    .QN_t(n6121_t)
  );


  sdffs1
  \DFF_217/Q_reg 
  (
    .DIN(WX1827),
    .DIN_t(WX1827_t),
    .SDIN(n6995),
    .SDIN_t(n6995_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6996),
    .Q_t(n6996_t),
    .QN(n6122),
    .QN_t(n6122_t)
  );


  sdffs1
  \DFF_216/Q_reg 
  (
    .DIN(WX1825),
    .DIN_t(WX1825_t),
    .SDIN(n6994),
    .SDIN_t(n6994_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6995),
    .Q_t(n6995_t),
    .QN(n6123),
    .QN_t(n6123_t)
  );


  sdffs1
  \DFF_215/Q_reg 
  (
    .DIN(WX1823),
    .DIN_t(WX1823_t),
    .SDIN(n6993),
    .SDIN_t(n6993_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6994),
    .Q_t(n6994_t),
    .QN(n6124),
    .QN_t(n6124_t)
  );


  sdffs1
  \DFF_214/Q_reg 
  (
    .DIN(WX1821),
    .DIN_t(WX1821_t),
    .SDIN(n6992),
    .SDIN_t(n6992_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6993),
    .Q_t(n6993_t),
    .QN(n6125),
    .QN_t(n6125_t)
  );


  sdffs1
  \DFF_213/Q_reg 
  (
    .DIN(WX1819),
    .DIN_t(WX1819_t),
    .SDIN(n6991),
    .SDIN_t(n6991_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6992),
    .Q_t(n6992_t),
    .QN(n6126),
    .QN_t(n6126_t)
  );


  sdffs1
  \DFF_212/Q_reg 
  (
    .DIN(WX1817),
    .DIN_t(WX1817_t),
    .SDIN(n6990),
    .SDIN_t(n6990_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6991),
    .Q_t(n6991_t),
    .QN(n6127),
    .QN_t(n6127_t)
  );


  sdffs1
  \DFF_211/Q_reg 
  (
    .DIN(WX1815),
    .DIN_t(WX1815_t),
    .SDIN(n6989),
    .SDIN_t(n6989_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6990),
    .Q_t(n6990_t),
    .QN(n6128),
    .QN_t(n6128_t)
  );


  sdffs1
  \DFF_210/Q_reg 
  (
    .DIN(WX1813),
    .DIN_t(WX1813_t),
    .SDIN(n6988),
    .SDIN_t(n6988_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6989),
    .Q_t(n6989_t),
    .QN(n6129),
    .QN_t(n6129_t)
  );


  sdffs1
  \DFF_209/Q_reg 
  (
    .DIN(WX1811),
    .DIN_t(WX1811_t),
    .SDIN(n6987),
    .SDIN_t(n6987_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6988),
    .Q_t(n6988_t),
    .QN(n6130),
    .QN_t(n6130_t)
  );


  sdffs1
  \DFF_208/Q_reg 
  (
    .DIN(WX1809),
    .DIN_t(WX1809_t),
    .SDIN(n6986),
    .SDIN_t(n6986_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6987),
    .Q_t(n6987_t),
    .QN(n6131),
    .QN_t(n6131_t)
  );


  sdffs1
  \DFF_207/Q_reg 
  (
    .DIN(WX1807),
    .DIN_t(WX1807_t),
    .SDIN(n6985),
    .SDIN_t(n6985_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6986),
    .Q_t(n6986_t),
    .QN(n6132),
    .QN_t(n6132_t)
  );


  sdffs1
  \DFF_206/Q_reg 
  (
    .DIN(WX1805),
    .DIN_t(WX1805_t),
    .SDIN(n6984),
    .SDIN_t(n6984_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6985),
    .Q_t(n6985_t),
    .QN(n6133),
    .QN_t(n6133_t)
  );


  sdffs1
  \DFF_205/Q_reg 
  (
    .DIN(WX1803),
    .DIN_t(WX1803_t),
    .SDIN(n6983),
    .SDIN_t(n6983_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6984),
    .Q_t(n6984_t),
    .QN(n6134),
    .QN_t(n6134_t)
  );


  sdffs1
  \DFF_204/Q_reg 
  (
    .DIN(WX1801),
    .DIN_t(WX1801_t),
    .SDIN(n6982),
    .SDIN_t(n6982_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6983),
    .Q_t(n6983_t),
    .QN(n6135),
    .QN_t(n6135_t)
  );


  sdffs1
  \DFF_203/Q_reg 
  (
    .DIN(WX1799),
    .DIN_t(WX1799_t),
    .SDIN(n6981),
    .SDIN_t(n6981_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6982),
    .Q_t(n6982_t),
    .QN(n6136),
    .QN_t(n6136_t)
  );


  sdffs1
  \DFF_202/Q_reg 
  (
    .DIN(WX1797),
    .DIN_t(WX1797_t),
    .SDIN(n6980),
    .SDIN_t(n6980_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6981),
    .Q_t(n6981_t),
    .QN(n6137),
    .QN_t(n6137_t)
  );


  sdffs1
  \DFF_201/Q_reg 
  (
    .DIN(WX1795),
    .DIN_t(WX1795_t),
    .SDIN(n6979),
    .SDIN_t(n6979_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6980),
    .Q_t(n6980_t),
    .QN(n6138),
    .QN_t(n6138_t)
  );


  sdffs1
  \DFF_200/Q_reg 
  (
    .DIN(WX1793),
    .DIN_t(WX1793_t),
    .SDIN(n6978),
    .SDIN_t(n6978_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6979),
    .Q_t(n6979_t),
    .QN(n6139),
    .QN_t(n6139_t)
  );


  sdffs1
  \DFF_199/Q_reg 
  (
    .DIN(WX1791),
    .DIN_t(WX1791_t),
    .SDIN(n6977),
    .SDIN_t(n6977_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6978),
    .Q_t(n6978_t),
    .QN(n6140),
    .QN_t(n6140_t)
  );


  sdffs1
  \DFF_198/Q_reg 
  (
    .DIN(WX1789),
    .DIN_t(WX1789_t),
    .SDIN(n6976),
    .SDIN_t(n6976_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6977),
    .Q_t(n6977_t),
    .QN(n6141),
    .QN_t(n6141_t)
  );


  sdffs1
  \DFF_197/Q_reg 
  (
    .DIN(WX1787),
    .DIN_t(WX1787_t),
    .SDIN(n6975),
    .SDIN_t(n6975_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6976),
    .Q_t(n6976_t),
    .QN(n6142),
    .QN_t(n6142_t)
  );


  sdffs1
  \DFF_196/Q_reg 
  (
    .DIN(WX1785),
    .DIN_t(WX1785_t),
    .SDIN(n6974),
    .SDIN_t(n6974_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6975),
    .Q_t(n6975_t),
    .QN(n6143),
    .QN_t(n6143_t)
  );


  sdffs1
  \DFF_195/Q_reg 
  (
    .DIN(WX1783),
    .DIN_t(WX1783_t),
    .SDIN(n6973),
    .SDIN_t(n6973_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6974),
    .Q_t(n6974_t),
    .QN(n6144),
    .QN_t(n6144_t)
  );


  sdffs1
  \DFF_194/Q_reg 
  (
    .DIN(WX1781),
    .DIN_t(WX1781_t),
    .SDIN(n6972),
    .SDIN_t(n6972_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6973),
    .Q_t(n6973_t),
    .QN(n6145),
    .QN_t(n6145_t)
  );


  sdffs1
  \DFF_193/Q_reg 
  (
    .DIN(WX1779),
    .DIN_t(WX1779_t),
    .SDIN(n6971),
    .SDIN_t(n6971_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6972),
    .Q_t(n6972_t),
    .QN(n6146),
    .QN_t(n6146_t)
  );


  sdffs1
  \DFF_192/Q_reg 
  (
    .DIN(WX1777),
    .DIN_t(WX1777_t),
    .SDIN(CRC_OUT_9_31),
    .SDIN_t(CRC_OUT_9_31_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6971),
    .Q_t(n6971_t),
    .QN(n6115),
    .QN_t(n6115_t)
  );


  sdffs1
  \DFF_191/Q_reg 
  (
    .DIN(WX1326),
    .DIN_t(WX1326_t),
    .SDIN(CRC_OUT_9_30),
    .SDIN_t(CRC_OUT_9_30_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_31),
    .Q_t(CRC_OUT_9_31_t),
    .QN(n6178),
    .QN_t(n6178_t)
  );


  sdffs1
  \DFF_190/Q_reg 
  (
    .DIN(WX1324),
    .DIN_t(WX1324_t),
    .SDIN(CRC_OUT_9_29),
    .SDIN_t(CRC_OUT_9_29_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_30),
    .Q_t(CRC_OUT_9_30_t),
    .QN(n6147),
    .QN_t(n6147_t)
  );


  sdffs1
  \DFF_189/Q_reg 
  (
    .DIN(WX1322),
    .DIN_t(WX1322_t),
    .SDIN(CRC_OUT_9_28),
    .SDIN_t(CRC_OUT_9_28_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_29),
    .Q_t(CRC_OUT_9_29_t),
    .QN(n6148),
    .QN_t(n6148_t)
  );


  sdffs1
  \DFF_188/Q_reg 
  (
    .DIN(WX1320),
    .DIN_t(WX1320_t),
    .SDIN(CRC_OUT_9_27),
    .SDIN_t(CRC_OUT_9_27_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_28),
    .Q_t(CRC_OUT_9_28_t),
    .QN(n6149),
    .QN_t(n6149_t)
  );


  sdffs1
  \DFF_187/Q_reg 
  (
    .DIN(WX1318),
    .DIN_t(WX1318_t),
    .SDIN(CRC_OUT_9_26),
    .SDIN_t(CRC_OUT_9_26_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_27),
    .Q_t(CRC_OUT_9_27_t),
    .QN(n6150),
    .QN_t(n6150_t)
  );


  sdffs1
  \DFF_186/Q_reg 
  (
    .DIN(WX1316),
    .DIN_t(WX1316_t),
    .SDIN(CRC_OUT_9_25),
    .SDIN_t(CRC_OUT_9_25_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_26),
    .Q_t(CRC_OUT_9_26_t),
    .QN(n6151),
    .QN_t(n6151_t)
  );


  sdffs1
  \DFF_185/Q_reg 
  (
    .DIN(WX1314),
    .DIN_t(WX1314_t),
    .SDIN(CRC_OUT_9_24),
    .SDIN_t(CRC_OUT_9_24_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_25),
    .Q_t(CRC_OUT_9_25_t),
    .QN(n6152),
    .QN_t(n6152_t)
  );


  sdffs1
  \DFF_184/Q_reg 
  (
    .DIN(WX1312),
    .DIN_t(WX1312_t),
    .SDIN(CRC_OUT_9_23),
    .SDIN_t(CRC_OUT_9_23_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_24),
    .Q_t(CRC_OUT_9_24_t),
    .QN(n6153),
    .QN_t(n6153_t)
  );


  sdffs1
  \DFF_183/Q_reg 
  (
    .DIN(WX1310),
    .DIN_t(WX1310_t),
    .SDIN(CRC_OUT_9_22),
    .SDIN_t(CRC_OUT_9_22_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_23),
    .Q_t(CRC_OUT_9_23_t),
    .QN(n6154),
    .QN_t(n6154_t)
  );


  sdffs1
  \DFF_182/Q_reg 
  (
    .DIN(WX1308),
    .DIN_t(WX1308_t),
    .SDIN(CRC_OUT_9_21),
    .SDIN_t(CRC_OUT_9_21_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_22),
    .Q_t(CRC_OUT_9_22_t),
    .QN(n6155),
    .QN_t(n6155_t)
  );


  sdffs1
  \DFF_181/Q_reg 
  (
    .DIN(WX1306),
    .DIN_t(WX1306_t),
    .SDIN(CRC_OUT_9_20),
    .SDIN_t(CRC_OUT_9_20_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_21),
    .Q_t(CRC_OUT_9_21_t),
    .QN(n6156),
    .QN_t(n6156_t)
  );


  sdffs1
  \DFF_180/Q_reg 
  (
    .DIN(WX1304),
    .DIN_t(WX1304_t),
    .SDIN(CRC_OUT_9_19),
    .SDIN_t(CRC_OUT_9_19_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_20),
    .Q_t(CRC_OUT_9_20_t),
    .QN(n6157),
    .QN_t(n6157_t)
  );


  sdffs1
  \DFF_179/Q_reg 
  (
    .DIN(WX1302),
    .DIN_t(WX1302_t),
    .SDIN(CRC_OUT_9_18),
    .SDIN_t(CRC_OUT_9_18_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_19),
    .Q_t(CRC_OUT_9_19_t),
    .QN(n6158),
    .QN_t(n6158_t)
  );


  sdffs1
  \DFF_178/Q_reg 
  (
    .DIN(WX1300),
    .DIN_t(WX1300_t),
    .SDIN(CRC_OUT_9_17),
    .SDIN_t(CRC_OUT_9_17_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_18),
    .Q_t(CRC_OUT_9_18_t),
    .QN(n6159),
    .QN_t(n6159_t)
  );


  sdffs1
  \DFF_177/Q_reg 
  (
    .DIN(WX1298),
    .DIN_t(WX1298_t),
    .SDIN(CRC_OUT_9_16),
    .SDIN_t(CRC_OUT_9_16_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_17),
    .Q_t(CRC_OUT_9_17_t),
    .QN(n6160),
    .QN_t(n6160_t)
  );


  sdffs1
  \DFF_176/Q_reg 
  (
    .DIN(WX1296),
    .DIN_t(WX1296_t),
    .SDIN(CRC_OUT_9_15),
    .SDIN_t(CRC_OUT_9_15_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_16),
    .Q_t(CRC_OUT_9_16_t),
    .QN(n6161),
    .QN_t(n6161_t)
  );


  sdffs1
  \DFF_175/Q_reg 
  (
    .DIN(WX1294),
    .DIN_t(WX1294_t),
    .SDIN(CRC_OUT_9_14),
    .SDIN_t(CRC_OUT_9_14_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_15),
    .Q_t(CRC_OUT_9_15_t),
    .QN(n6162),
    .QN_t(n6162_t)
  );


  sdffs1
  \DFF_174/Q_reg 
  (
    .DIN(WX1292),
    .DIN_t(WX1292_t),
    .SDIN(CRC_OUT_9_13),
    .SDIN_t(CRC_OUT_9_13_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_14),
    .Q_t(CRC_OUT_9_14_t),
    .QN(n6163),
    .QN_t(n6163_t)
  );


  sdffs1
  \DFF_173/Q_reg 
  (
    .DIN(WX1290),
    .DIN_t(WX1290_t),
    .SDIN(CRC_OUT_9_12),
    .SDIN_t(CRC_OUT_9_12_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_13),
    .Q_t(CRC_OUT_9_13_t),
    .QN(n6164),
    .QN_t(n6164_t)
  );


  sdffs1
  \DFF_172/Q_reg 
  (
    .DIN(WX1288),
    .DIN_t(WX1288_t),
    .SDIN(CRC_OUT_9_11),
    .SDIN_t(CRC_OUT_9_11_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_12),
    .Q_t(CRC_OUT_9_12_t),
    .QN(n6165),
    .QN_t(n6165_t)
  );


  sdffs1
  \DFF_171/Q_reg 
  (
    .DIN(WX1286),
    .DIN_t(WX1286_t),
    .SDIN(CRC_OUT_9_10),
    .SDIN_t(CRC_OUT_9_10_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_11),
    .Q_t(CRC_OUT_9_11_t),
    .QN(n6166),
    .QN_t(n6166_t)
  );


  sdffs1
  \DFF_170/Q_reg 
  (
    .DIN(WX1284),
    .DIN_t(WX1284_t),
    .SDIN(CRC_OUT_9_9),
    .SDIN_t(CRC_OUT_9_9_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_10),
    .Q_t(CRC_OUT_9_10_t),
    .QN(n6167),
    .QN_t(n6167_t)
  );


  sdffs1
  \DFF_169/Q_reg 
  (
    .DIN(WX1282),
    .DIN_t(WX1282_t),
    .SDIN(CRC_OUT_9_8),
    .SDIN_t(CRC_OUT_9_8_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_9),
    .Q_t(CRC_OUT_9_9_t),
    .QN(n6168),
    .QN_t(n6168_t)
  );


  sdffs1
  \DFF_168/Q_reg 
  (
    .DIN(WX1280),
    .DIN_t(WX1280_t),
    .SDIN(CRC_OUT_9_7),
    .SDIN_t(CRC_OUT_9_7_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_8),
    .Q_t(CRC_OUT_9_8_t),
    .QN(n6169),
    .QN_t(n6169_t)
  );


  sdffs1
  \DFF_167/Q_reg 
  (
    .DIN(WX1278),
    .DIN_t(WX1278_t),
    .SDIN(CRC_OUT_9_6),
    .SDIN_t(CRC_OUT_9_6_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_7),
    .Q_t(CRC_OUT_9_7_t),
    .QN(n6170),
    .QN_t(n6170_t)
  );


  sdffs1
  \DFF_166/Q_reg 
  (
    .DIN(WX1276),
    .DIN_t(WX1276_t),
    .SDIN(CRC_OUT_9_5),
    .SDIN_t(CRC_OUT_9_5_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_6),
    .Q_t(CRC_OUT_9_6_t),
    .QN(n6171),
    .QN_t(n6171_t)
  );


  sdffs1
  \DFF_165/Q_reg 
  (
    .DIN(WX1274),
    .DIN_t(WX1274_t),
    .SDIN(CRC_OUT_9_4),
    .SDIN_t(CRC_OUT_9_4_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_5),
    .Q_t(CRC_OUT_9_5_t),
    .QN(n6172),
    .QN_t(n6172_t)
  );


  sdffs1
  \DFF_164/Q_reg 
  (
    .DIN(WX1272),
    .DIN_t(WX1272_t),
    .SDIN(CRC_OUT_9_3),
    .SDIN_t(CRC_OUT_9_3_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_4),
    .Q_t(CRC_OUT_9_4_t),
    .QN(n6173),
    .QN_t(n6173_t)
  );


  sdffs1
  \DFF_163/Q_reg 
  (
    .DIN(WX1270),
    .DIN_t(WX1270_t),
    .SDIN(CRC_OUT_9_2),
    .SDIN_t(CRC_OUT_9_2_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_3),
    .Q_t(CRC_OUT_9_3_t),
    .QN(n6174),
    .QN_t(n6174_t)
  );


  sdffs1
  \DFF_162/Q_reg 
  (
    .DIN(WX1268),
    .DIN_t(WX1268_t),
    .SDIN(CRC_OUT_9_1),
    .SDIN_t(CRC_OUT_9_1_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_2),
    .Q_t(CRC_OUT_9_2_t),
    .QN(n6175),
    .QN_t(n6175_t)
  );


  sdffs1
  \DFF_161/Q_reg 
  (
    .DIN(WX1266),
    .DIN_t(WX1266_t),
    .SDIN(CRC_OUT_9_0),
    .SDIN_t(CRC_OUT_9_0_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_1),
    .Q_t(CRC_OUT_9_1_t),
    .QN(n6176),
    .QN_t(n6176_t)
  );


  sdffs1
  \DFF_160/Q_reg 
  (
    .DIN(WX1264),
    .DIN_t(WX1264_t),
    .SDIN(n6970),
    .SDIN_t(n6970_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(CRC_OUT_9_0),
    .Q_t(CRC_OUT_9_0_t),
    .QN(n6177),
    .QN_t(n6177_t)
  );


  sdffs1
  \DFF_159/Q_reg 
  (
    .DIN(WX898),
    .DIN_t(WX898_t),
    .SDIN(n6969),
    .SDIN_t(n6969_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6970),
    .Q_t(n6970_t),
    .QN(n6462),
    .QN_t(n6462_t)
  );


  sdffs1
  \DFF_158/Q_reg 
  (
    .DIN(WX896),
    .DIN_t(WX896_t),
    .SDIN(n6968),
    .SDIN_t(n6968_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6969),
    .Q_t(n6969_t),
    .QN(n6530),
    .QN_t(n6530_t)
  );


  sdffs1
  \DFF_157/Q_reg 
  (
    .DIN(WX894),
    .DIN_t(WX894_t),
    .SDIN(n6967),
    .SDIN_t(n6967_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6968),
    .Q_t(n6968_t),
    .QN(n6437),
    .QN_t(n6437_t)
  );


  sdffs1
  \DFF_156/Q_reg 
  (
    .DIN(WX892),
    .DIN_t(WX892_t),
    .SDIN(n6966),
    .SDIN_t(n6966_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6967),
    .Q_t(n6967_t),
    .QN(n6468),
    .QN_t(n6468_t)
  );


  sdffs1
  \DFF_155/Q_reg 
  (
    .DIN(WX890),
    .DIN_t(WX890_t),
    .SDIN(n6965),
    .SDIN_t(n6965_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6966),
    .Q_t(n6966_t),
    .QN(n6471),
    .QN_t(n6471_t)
  );


  sdffs1
  \DFF_154/Q_reg 
  (
    .DIN(WX888),
    .DIN_t(WX888_t),
    .SDIN(n6964),
    .SDIN_t(n6964_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6965),
    .Q_t(n6965_t),
    .QN(n6459),
    .QN_t(n6459_t)
  );


  sdffs1
  \DFF_153/Q_reg 
  (
    .DIN(WX886),
    .DIN_t(WX886_t),
    .SDIN(n6963),
    .SDIN_t(n6963_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6964),
    .Q_t(n6964_t),
    .QN(n6441),
    .QN_t(n6441_t)
  );


  sdffs1
  \DFF_152/Q_reg 
  (
    .DIN(WX884),
    .DIN_t(WX884_t),
    .SDIN(n6962),
    .SDIN_t(n6962_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6963),
    .Q_t(n6963_t),
    .QN(n6465),
    .QN_t(n6465_t)
  );


  sdffs1
  \DFF_151/Q_reg 
  (
    .DIN(WX882),
    .DIN_t(WX882_t),
    .SDIN(n6961),
    .SDIN_t(n6961_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6962),
    .Q_t(n6962_t),
    .QN(n6453),
    .QN_t(n6453_t)
  );


  sdffs1
  \DFF_150/Q_reg 
  (
    .DIN(WX880),
    .DIN_t(WX880_t),
    .SDIN(n6960),
    .SDIN_t(n6960_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6961),
    .Q_t(n6961_t),
    .QN(n6506),
    .QN_t(n6506_t)
  );


  sdffs1
  \DFF_149/Q_reg 
  (
    .DIN(WX878),
    .DIN_t(WX878_t),
    .SDIN(n6959),
    .SDIN_t(n6959_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6960),
    .Q_t(n6960_t),
    .QN(n6450),
    .QN_t(n6450_t)
  );


  sdffs1
  \DFF_148/Q_reg 
  (
    .DIN(WX876),
    .DIN_t(WX876_t),
    .SDIN(n6958),
    .SDIN_t(n6958_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6959),
    .Q_t(n6959_t),
    .QN(n6444),
    .QN_t(n6444_t)
  );


  sdffs1
  \DFF_147/Q_reg 
  (
    .DIN(WX874),
    .DIN_t(WX874_t),
    .SDIN(n6957),
    .SDIN_t(n6957_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6958),
    .Q_t(n6958_t),
    .QN(n6456),
    .QN_t(n6456_t)
  );


  sdffs1
  \DFF_146/Q_reg 
  (
    .DIN(WX872),
    .DIN_t(WX872_t),
    .SDIN(n6956),
    .SDIN_t(n6956_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6957),
    .Q_t(n6957_t),
    .QN(n6447),
    .QN_t(n6447_t)
  );


  sdffs1
  \DFF_145/Q_reg 
  (
    .DIN(WX870),
    .DIN_t(WX870_t),
    .SDIN(n6955),
    .SDIN_t(n6955_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6956),
    .Q_t(n6956_t),
    .QN(n6525),
    .QN_t(n6525_t)
  );


  sdffs1
  \DFF_144/Q_reg 
  (
    .DIN(WX868),
    .DIN_t(WX868_t),
    .SDIN(n6954),
    .SDIN_t(n6954_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6955),
    .Q_t(n6955_t),
    .QN(n6438),
    .QN_t(n6438_t)
  );


  sdffs1
  \DFF_143/Q_reg 
  (
    .DIN(WX866),
    .DIN_t(WX866_t),
    .SDIN(n6953),
    .SDIN_t(n6953_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6954),
    .Q_t(n6954_t),
    .QN(n6510),
    .QN_t(n6510_t)
  );


  sdffs1
  \DFF_142/Q_reg 
  (
    .DIN(WX864),
    .DIN_t(WX864_t),
    .SDIN(n6952),
    .SDIN_t(n6952_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6953),
    .Q_t(n6953_t),
    .QN(n6495),
    .QN_t(n6495_t)
  );


  sdffs1
  \DFF_141/Q_reg 
  (
    .DIN(WX862),
    .DIN_t(WX862_t),
    .SDIN(n6951),
    .SDIN_t(n6951_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6952),
    .Q_t(n6952_t),
    .QN(n6491),
    .QN_t(n6491_t)
  );


  sdffs1
  \DFF_140/Q_reg 
  (
    .DIN(WX860),
    .DIN_t(WX860_t),
    .SDIN(n6950),
    .SDIN_t(n6950_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6951),
    .Q_t(n6951_t),
    .QN(n6477),
    .QN_t(n6477_t)
  );


  sdffs1
  \DFF_139/Q_reg 
  (
    .DIN(WX858),
    .DIN_t(WX858_t),
    .SDIN(n6949),
    .SDIN_t(n6949_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6950),
    .Q_t(n6950_t),
    .QN(n6522),
    .QN_t(n6522_t)
  );


  sdffs1
  \DFF_138/Q_reg 
  (
    .DIN(WX856),
    .DIN_t(WX856_t),
    .SDIN(n6948),
    .SDIN_t(n6948_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6949),
    .Q_t(n6949_t),
    .QN(n6517),
    .QN_t(n6517_t)
  );


  sdffs1
  \DFF_137/Q_reg 
  (
    .DIN(WX854),
    .DIN_t(WX854_t),
    .SDIN(n6947),
    .SDIN_t(n6947_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6948),
    .Q_t(n6948_t),
    .QN(n6516),
    .QN_t(n6516_t)
  );


  sdffs1
  \DFF_136/Q_reg 
  (
    .DIN(WX852),
    .DIN_t(WX852_t),
    .SDIN(n6946),
    .SDIN_t(n6946_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6947),
    .Q_t(n6947_t),
    .QN(n6511),
    .QN_t(n6511_t)
  );


  sdffs1
  \DFF_135/Q_reg 
  (
    .DIN(WX850),
    .DIN_t(WX850_t),
    .SDIN(n6945),
    .SDIN_t(n6945_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6946),
    .Q_t(n6946_t),
    .QN(n6501),
    .QN_t(n6501_t)
  );


  sdffs1
  \DFF_134/Q_reg 
  (
    .DIN(WX848),
    .DIN_t(WX848_t),
    .SDIN(n6944),
    .SDIN_t(n6944_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6945),
    .Q_t(n6945_t),
    .QN(n6500),
    .QN_t(n6500_t)
  );


  sdffs1
  \DFF_133/Q_reg 
  (
    .DIN(WX846),
    .DIN_t(WX846_t),
    .SDIN(n6943),
    .SDIN_t(n6943_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6944),
    .Q_t(n6944_t),
    .QN(n6492),
    .QN_t(n6492_t)
  );


  sdffs1
  \DFF_132/Q_reg 
  (
    .DIN(WX844),
    .DIN_t(WX844_t),
    .SDIN(n6942),
    .SDIN_t(n6942_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6943),
    .Q_t(n6943_t),
    .QN(n6486),
    .QN_t(n6486_t)
  );


  sdffs1
  \DFF_131/Q_reg 
  (
    .DIN(WX842),
    .DIN_t(WX842_t),
    .SDIN(n6941),
    .SDIN_t(n6941_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6942),
    .Q_t(n6942_t),
    .QN(n6483),
    .QN_t(n6483_t)
  );


  sdffs1
  \DFF_130/Q_reg 
  (
    .DIN(WX840),
    .DIN_t(WX840_t),
    .SDIN(n6940),
    .SDIN_t(n6940_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6941),
    .Q_t(n6941_t),
    .QN(n6482),
    .QN_t(n6482_t)
  );


  sdffs1
  \DFF_129/Q_reg 
  (
    .DIN(WX838),
    .DIN_t(WX838_t),
    .SDIN(n6939),
    .SDIN_t(n6939_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6940),
    .Q_t(n6940_t),
    .QN(n6474),
    .QN_t(n6474_t)
  );


  sdffs1
  \DFF_128/Q_reg 
  (
    .DIN(WX836),
    .DIN_t(WX836_t),
    .SDIN(n6938),
    .SDIN_t(n6938_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6939),
    .Q_t(n6939_t),
    .QN(n6534),
    .QN_t(n6534_t)
  );


  sdffs1
  \DFF_127/Q_reg 
  (
    .DIN(WX834),
    .DIN_t(WX834_t),
    .SDIN(n6937),
    .SDIN_t(n6937_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6938),
    .Q_t(n6938_t),
    .QN(n6463),
    .QN_t(n6463_t)
  );


  sdffs1
  \DFF_126/Q_reg 
  (
    .DIN(WX832),
    .DIN_t(WX832_t),
    .SDIN(n6936),
    .SDIN_t(n6936_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6937),
    .Q_t(n6937_t),
    .QN(n6527),
    .QN_t(n6527_t)
  );


  sdffs1
  \DFF_125/Q_reg 
  (
    .DIN(WX830),
    .DIN_t(WX830_t),
    .SDIN(n6935),
    .SDIN_t(n6935_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6936),
    .Q_t(n6936_t),
    .QN(n6436),
    .QN_t(n6436_t)
  );


  sdffs1
  \DFF_124/Q_reg 
  (
    .DIN(WX828),
    .DIN_t(WX828_t),
    .SDIN(n6934),
    .SDIN_t(n6934_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6935),
    .Q_t(n6935_t),
    .QN(n6469),
    .QN_t(n6469_t)
  );


  sdffs1
  \DFF_123/Q_reg 
  (
    .DIN(WX826),
    .DIN_t(WX826_t),
    .SDIN(n6933),
    .SDIN_t(n6933_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6934),
    .Q_t(n6934_t),
    .QN(n6472),
    .QN_t(n6472_t)
  );


  sdffs1
  \DFF_122/Q_reg 
  (
    .DIN(WX824),
    .DIN_t(WX824_t),
    .SDIN(n6932),
    .SDIN_t(n6932_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6933),
    .Q_t(n6933_t),
    .QN(n6460),
    .QN_t(n6460_t)
  );


  sdffs1
  \DFF_121/Q_reg 
  (
    .DIN(WX822),
    .DIN_t(WX822_t),
    .SDIN(n6931),
    .SDIN_t(n6931_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6932),
    .Q_t(n6932_t),
    .QN(n6442),
    .QN_t(n6442_t)
  );


  sdffs1
  \DFF_120/Q_reg 
  (
    .DIN(WX820),
    .DIN_t(WX820_t),
    .SDIN(n6930),
    .SDIN_t(n6930_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6931),
    .Q_t(n6931_t),
    .QN(n6466),
    .QN_t(n6466_t)
  );


  sdffs1
  \DFF_119/Q_reg 
  (
    .DIN(WX818),
    .DIN_t(WX818_t),
    .SDIN(n6929),
    .SDIN_t(n6929_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6930),
    .Q_t(n6930_t),
    .QN(n6454),
    .QN_t(n6454_t)
  );


  sdffs1
  \DFF_118/Q_reg 
  (
    .DIN(WX816),
    .DIN_t(WX816_t),
    .SDIN(n6928),
    .SDIN_t(n6928_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6929),
    .Q_t(n6929_t),
    .QN(n6504),
    .QN_t(n6504_t)
  );


  sdffs1
  \DFF_117/Q_reg 
  (
    .DIN(WX814),
    .DIN_t(WX814_t),
    .SDIN(n6927),
    .SDIN_t(n6927_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6928),
    .Q_t(n6928_t),
    .QN(n6451),
    .QN_t(n6451_t)
  );


  sdffs1
  \DFF_116/Q_reg 
  (
    .DIN(WX812),
    .DIN_t(WX812_t),
    .SDIN(n6926),
    .SDIN_t(n6926_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6927),
    .Q_t(n6927_t),
    .QN(n6445),
    .QN_t(n6445_t)
  );


  sdffs1
  \DFF_115/Q_reg 
  (
    .DIN(WX810),
    .DIN_t(WX810_t),
    .SDIN(n6925),
    .SDIN_t(n6925_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6926),
    .Q_t(n6926_t),
    .QN(n6457),
    .QN_t(n6457_t)
  );


  sdffs1
  \DFF_114/Q_reg 
  (
    .DIN(WX808),
    .DIN_t(WX808_t),
    .SDIN(n6924),
    .SDIN_t(n6924_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6925),
    .Q_t(n6925_t),
    .QN(n6448),
    .QN_t(n6448_t)
  );


  sdffs1
  \DFF_113/Q_reg 
  (
    .DIN(WX806),
    .DIN_t(WX806_t),
    .SDIN(n6923),
    .SDIN_t(n6923_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6924),
    .Q_t(n6924_t),
    .QN(n6523),
    .QN_t(n6523_t)
  );


  sdffs1
  \DFF_112/Q_reg 
  (
    .DIN(WX804),
    .DIN_t(WX804_t),
    .SDIN(n6922),
    .SDIN_t(n6922_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6923),
    .Q_t(n6923_t),
    .QN(n6439),
    .QN_t(n6439_t)
  );


  sdffs1
  \DFF_111/Q_reg 
  (
    .DIN(WX802),
    .DIN_t(WX802_t),
    .SDIN(n6921),
    .SDIN_t(n6921_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6922),
    .Q_t(n6922_t),
    .QN(n6539),
    .QN_t(n6539_t)
  );


  sdffs1
  \DFF_110/Q_reg 
  (
    .DIN(WX800),
    .DIN_t(WX800_t),
    .SDIN(n6920),
    .SDIN_t(n6920_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6921),
    .Q_t(n6921_t),
    .QN(n6496),
    .QN_t(n6496_t)
  );


  sdffs1
  \DFF_109/Q_reg 
  (
    .DIN(WX798),
    .DIN_t(WX798_t),
    .SDIN(n6919),
    .SDIN_t(n6919_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6920),
    .Q_t(n6920_t),
    .QN(n6544),
    .QN_t(n6544_t)
  );


  sdffs1
  \DFF_108/Q_reg 
  (
    .DIN(WX796),
    .DIN_t(WX796_t),
    .SDIN(n6918),
    .SDIN_t(n6918_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6919),
    .Q_t(n6919_t),
    .QN(n6478),
    .QN_t(n6478_t)
  );


  sdffs1
  \DFF_107/Q_reg 
  (
    .DIN(WX794),
    .DIN_t(WX794_t),
    .SDIN(n6917),
    .SDIN_t(n6917_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6918),
    .Q_t(n6918_t),
    .QN(n6535),
    .QN_t(n6535_t)
  );


  sdffs1
  \DFF_106/Q_reg 
  (
    .DIN(WX792),
    .DIN_t(WX792_t),
    .SDIN(n6916),
    .SDIN_t(n6916_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6917),
    .Q_t(n6917_t),
    .QN(n6518),
    .QN_t(n6518_t)
  );


  sdffs1
  \DFF_105/Q_reg 
  (
    .DIN(WX790),
    .DIN_t(WX790_t),
    .SDIN(n6915),
    .SDIN_t(n6915_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6916),
    .Q_t(n6916_t),
    .QN(n6537),
    .QN_t(n6537_t)
  );


  sdffs1
  \DFF_104/Q_reg 
  (
    .DIN(WX788),
    .DIN_t(WX788_t),
    .SDIN(n6914),
    .SDIN_t(n6914_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6915),
    .Q_t(n6915_t),
    .QN(n6512),
    .QN_t(n6512_t)
  );


  sdffs1
  \DFF_103/Q_reg 
  (
    .DIN(WX786),
    .DIN_t(WX786_t),
    .SDIN(n6913),
    .SDIN_t(n6913_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6914),
    .Q_t(n6914_t),
    .QN(n6502),
    .QN_t(n6502_t)
  );


  sdffs1
  \DFF_102/Q_reg 
  (
    .DIN(WX784),
    .DIN_t(WX784_t),
    .SDIN(n6912),
    .SDIN_t(n6912_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6913),
    .Q_t(n6913_t),
    .QN(n6541),
    .QN_t(n6541_t)
  );


  sdffs1
  \DFF_101/Q_reg 
  (
    .DIN(WX782),
    .DIN_t(WX782_t),
    .SDIN(n6911),
    .SDIN_t(n6911_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6912),
    .Q_t(n6912_t),
    .QN(n6493),
    .QN_t(n6493_t)
  );


  sdffs1
  \DFF_100/Q_reg 
  (
    .DIN(WX780),
    .DIN_t(WX780_t),
    .SDIN(n6910),
    .SDIN_t(n6910_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6911),
    .Q_t(n6911_t),
    .QN(n6487),
    .QN_t(n6487_t)
  );


  sdffs1
  \DFF_99/Q_reg 
  (
    .DIN(WX778),
    .DIN_t(WX778_t),
    .SDIN(n6909),
    .SDIN_t(n6909_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6910),
    .Q_t(n6910_t),
    .QN(n6484),
    .QN_t(n6484_t)
  );


  sdffs1
  \DFF_98/Q_reg 
  (
    .DIN(WX776),
    .DIN_t(WX776_t),
    .SDIN(n6908),
    .SDIN_t(n6908_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6909),
    .Q_t(n6909_t),
    .QN(n6547),
    .QN_t(n6547_t)
  );


  sdffs1
  \DFF_97/Q_reg 
  (
    .DIN(WX774),
    .DIN_t(WX774_t),
    .SDIN(n6907),
    .SDIN_t(n6907_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6908),
    .Q_t(n6908_t),
    .QN(n6475),
    .QN_t(n6475_t)
  );


  sdffs1
  \DFF_96/Q_reg 
  (
    .DIN(WX772),
    .DIN_t(WX772_t),
    .SDIN(n6906),
    .SDIN_t(n6906_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6907),
    .Q_t(n6907_t),
    .QN(n6531),
    .QN_t(n6531_t)
  );


  sdffs1
  \DFF_95/Q_reg 
  (
    .DIN(WX770),
    .DIN_t(WX770_t),
    .SDIN(n6905),
    .SDIN_t(n6905_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6906),
    .Q_t(n6906_t),
    .QN(n6464),
    .QN_t(n6464_t)
  );


  sdffs1
  \DFF_94/Q_reg 
  (
    .DIN(WX768),
    .DIN_t(WX768_t),
    .SDIN(n6904),
    .SDIN_t(n6904_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6905),
    .Q_t(n6905_t),
    .QN(n6528),
    .QN_t(n6528_t)
  );


  sdffs1
  \DFF_93/Q_reg 
  (
    .DIN(WX766),
    .DIN_t(WX766_t),
    .SDIN(n6903),
    .SDIN_t(n6903_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6904),
    .Q_t(n6904_t),
    .QN(n6562),
    .QN_t(n6562_t)
  );


  sdffs1
  \DFF_92/Q_reg 
  (
    .DIN(WX764),
    .DIN_t(WX764_t),
    .SDIN(n6902),
    .SDIN_t(n6902_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6903),
    .Q_t(n6903_t),
    .QN(n6470),
    .QN_t(n6470_t)
  );


  sdffs1
  \DFF_91/Q_reg 
  (
    .DIN(WX762),
    .DIN_t(WX762_t),
    .SDIN(n6901),
    .SDIN_t(n6901_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6902),
    .Q_t(n6902_t),
    .QN(n6473),
    .QN_t(n6473_t)
  );


  sdffs1
  \DFF_90/Q_reg 
  (
    .DIN(WX760),
    .DIN_t(WX760_t),
    .SDIN(n6900),
    .SDIN_t(n6900_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6901),
    .Q_t(n6901_t),
    .QN(n6461),
    .QN_t(n6461_t)
  );


  sdffs1
  \DFF_89/Q_reg 
  (
    .DIN(WX758),
    .DIN_t(WX758_t),
    .SDIN(n6899),
    .SDIN_t(n6899_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6900),
    .Q_t(n6900_t),
    .QN(n6443),
    .QN_t(n6443_t)
  );


  sdffs1
  \DFF_88/Q_reg 
  (
    .DIN(WX756),
    .DIN_t(WX756_t),
    .SDIN(n6898),
    .SDIN_t(n6898_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6899),
    .Q_t(n6899_t),
    .QN(n6467),
    .QN_t(n6467_t)
  );


  sdffs1
  \DFF_87/Q_reg 
  (
    .DIN(WX754),
    .DIN_t(WX754_t),
    .SDIN(n6897),
    .SDIN_t(n6897_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6898),
    .Q_t(n6898_t),
    .QN(n6455),
    .QN_t(n6455_t)
  );


  sdffs1
  \DFF_86/Q_reg 
  (
    .DIN(WX752),
    .DIN_t(WX752_t),
    .SDIN(n6896),
    .SDIN_t(n6896_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6897),
    .Q_t(n6897_t),
    .QN(n6505),
    .QN_t(n6505_t)
  );


  sdffs1
  \DFF_85/Q_reg 
  (
    .DIN(WX750),
    .DIN_t(WX750_t),
    .SDIN(n6895),
    .SDIN_t(n6895_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6896),
    .Q_t(n6896_t),
    .QN(n6452),
    .QN_t(n6452_t)
  );


  sdffs1
  \DFF_84/Q_reg 
  (
    .DIN(WX748),
    .DIN_t(WX748_t),
    .SDIN(n6894),
    .SDIN_t(n6894_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6895),
    .Q_t(n6895_t),
    .QN(n6446),
    .QN_t(n6446_t)
  );


  sdffs1
  \DFF_83/Q_reg 
  (
    .DIN(WX746),
    .DIN_t(WX746_t),
    .SDIN(n6893),
    .SDIN_t(n6893_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6894),
    .Q_t(n6894_t),
    .QN(n6458),
    .QN_t(n6458_t)
  );


  sdffs1
  \DFF_82/Q_reg 
  (
    .DIN(WX744),
    .DIN_t(WX744_t),
    .SDIN(n6892),
    .SDIN_t(n6892_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6893),
    .Q_t(n6893_t),
    .QN(n6449),
    .QN_t(n6449_t)
  );


  sdffs1
  \DFF_81/Q_reg 
  (
    .DIN(WX742),
    .DIN_t(WX742_t),
    .SDIN(n6891),
    .SDIN_t(n6891_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6892),
    .Q_t(n6892_t),
    .QN(n6524),
    .QN_t(n6524_t)
  );


  sdffs1
  \DFF_80/Q_reg 
  (
    .DIN(WX740),
    .DIN_t(WX740_t),
    .SDIN(n6890),
    .SDIN_t(n6890_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6891),
    .Q_t(n6891_t),
    .QN(n6440),
    .QN_t(n6440_t)
  );


  sdffs1
  \DFF_79/Q_reg 
  (
    .DIN(WX738),
    .DIN_t(WX738_t),
    .SDIN(n6889),
    .SDIN_t(n6889_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6890),
    .Q_t(n6890_t),
    .QN(n6508),
    .QN_t(n6508_t)
  );


  sdffs1
  \DFF_78/Q_reg 
  (
    .DIN(WX736),
    .DIN_t(WX736_t),
    .SDIN(n6888),
    .SDIN_t(n6888_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6889),
    .Q_t(n6889_t),
    .QN(n6497),
    .QN_t(n6497_t)
  );


  sdffs1
  \DFF_77/Q_reg 
  (
    .DIN(WX734),
    .DIN_t(WX734_t),
    .SDIN(n6887),
    .SDIN_t(n6887_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6888),
    .Q_t(n6888_t),
    .QN(n6489),
    .QN_t(n6489_t)
  );


  sdffs1
  \DFF_76/Q_reg 
  (
    .DIN(WX732),
    .DIN_t(WX732_t),
    .SDIN(n6886),
    .SDIN_t(n6886_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6887),
    .Q_t(n6887_t),
    .QN(n6479),
    .QN_t(n6479_t)
  );


  sdffs1
  \DFF_75/Q_reg 
  (
    .DIN(WX730),
    .DIN_t(WX730_t),
    .SDIN(n6885),
    .SDIN_t(n6885_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6886),
    .Q_t(n6886_t),
    .QN(n6520),
    .QN_t(n6520_t)
  );


  sdffs1
  \DFF_74/Q_reg 
  (
    .DIN(WX728),
    .DIN_t(WX728_t),
    .SDIN(n6884),
    .SDIN_t(n6884_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6885),
    .Q_t(n6885_t),
    .QN(n6519),
    .QN_t(n6519_t)
  );


  sdffs1
  \DFF_73/Q_reg 
  (
    .DIN(WX726),
    .DIN_t(WX726_t),
    .SDIN(n6883),
    .SDIN_t(n6883_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6884),
    .Q_t(n6884_t),
    .QN(n6514),
    .QN_t(n6514_t)
  );


  sdffs1
  \DFF_72/Q_reg 
  (
    .DIN(WX724),
    .DIN_t(WX724_t),
    .SDIN(n6882),
    .SDIN_t(n6882_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6883),
    .Q_t(n6883_t),
    .QN(n6513),
    .QN_t(n6513_t)
  );


  sdffs1
  \DFF_71/Q_reg 
  (
    .DIN(WX722),
    .DIN_t(WX722_t),
    .SDIN(n6881),
    .SDIN_t(n6881_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6882),
    .Q_t(n6882_t),
    .QN(n6503),
    .QN_t(n6503_t)
  );


  sdffs1
  \DFF_70/Q_reg 
  (
    .DIN(WX720),
    .DIN_t(WX720_t),
    .SDIN(n6880),
    .SDIN_t(n6880_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6881),
    .Q_t(n6881_t),
    .QN(n6498),
    .QN_t(n6498_t)
  );


  sdffs1
  \DFF_69/Q_reg 
  (
    .DIN(WX718),
    .DIN_t(WX718_t),
    .SDIN(n6879),
    .SDIN_t(n6879_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6880),
    .Q_t(n6880_t),
    .QN(n6494),
    .QN_t(n6494_t)
  );


  sdffs1
  \DFF_68/Q_reg 
  (
    .DIN(WX716),
    .DIN_t(WX716_t),
    .SDIN(n6878),
    .SDIN_t(n6878_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6879),
    .Q_t(n6879_t),
    .QN(n6488),
    .QN_t(n6488_t)
  );


  sdffs1
  \DFF_67/Q_reg 
  (
    .DIN(WX714),
    .DIN_t(WX714_t),
    .SDIN(n6877),
    .SDIN_t(n6877_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6878),
    .Q_t(n6878_t),
    .QN(n6485),
    .QN_t(n6485_t)
  );


  sdffs1
  \DFF_66/Q_reg 
  (
    .DIN(WX712),
    .DIN_t(WX712_t),
    .SDIN(n6876),
    .SDIN_t(n6876_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6877),
    .Q_t(n6877_t),
    .QN(n6480),
    .QN_t(n6480_t)
  );


  sdffs1
  \DFF_65/Q_reg 
  (
    .DIN(WX710),
    .DIN_t(WX710_t),
    .SDIN(n6875),
    .SDIN_t(n6875_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6876),
    .Q_t(n6876_t),
    .QN(n6476),
    .QN_t(n6476_t)
  );


  sdffs1
  \DFF_64/Q_reg 
  (
    .DIN(WX708),
    .DIN_t(WX708_t),
    .SDIN(n6874),
    .SDIN_t(n6874_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6875),
    .Q_t(n6875_t),
    .QN(n6532),
    .QN_t(n6532_t)
  );


  sdffs1
  \DFF_63/Q_reg 
  (
    .DIN(WX706),
    .DIN_t(WX706_t),
    .SDIN(n6873),
    .SDIN_t(n6873_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6874),
    .Q_t(n6874_t),
    .QN(n6553),
    .QN_t(n6553_t)
  );


  sdffs1
  \DFF_62/Q_reg 
  (
    .DIN(WX704),
    .DIN_t(WX704_t),
    .SDIN(n6872),
    .SDIN_t(n6872_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6873),
    .Q_t(n6873_t),
    .QN(n6529),
    .QN_t(n6529_t)
  );


  sdffs1
  \DFF_61/Q_reg 
  (
    .DIN(WX702),
    .DIN_t(WX702_t),
    .SDIN(n6871),
    .SDIN_t(n6871_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6872),
    .Q_t(n6872_t),
    .QN(n6435),
    .QN_t(n6435_t)
  );


  sdffs1
  \DFF_60/Q_reg 
  (
    .DIN(WX700),
    .DIN_t(WX700_t),
    .SDIN(n6870),
    .SDIN_t(n6870_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6871),
    .Q_t(n6871_t),
    .QN(n6551),
    .QN_t(n6551_t)
  );


  sdffs1
  \DFF_59/Q_reg 
  (
    .DIN(WX698),
    .DIN_t(WX698_t),
    .SDIN(n6869),
    .SDIN_t(n6869_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6870),
    .Q_t(n6870_t),
    .QN(n6550),
    .QN_t(n6550_t)
  );


  sdffs1
  \DFF_58/Q_reg 
  (
    .DIN(WX696),
    .DIN_t(WX696_t),
    .SDIN(n6868),
    .SDIN_t(n6868_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6869),
    .Q_t(n6869_t),
    .QN(n6554),
    .QN_t(n6554_t)
  );


  sdffs1
  \DFF_57/Q_reg 
  (
    .DIN(WX694),
    .DIN_t(WX694_t),
    .SDIN(n6867),
    .SDIN_t(n6867_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6868),
    .Q_t(n6868_t),
    .QN(n6560),
    .QN_t(n6560_t)
  );


  sdffs1
  \DFF_56/Q_reg 
  (
    .DIN(WX692),
    .DIN_t(WX692_t),
    .SDIN(n6866),
    .SDIN_t(n6866_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6867),
    .Q_t(n6867_t),
    .QN(n6552),
    .QN_t(n6552_t)
  );


  sdffs1
  \DFF_55/Q_reg 
  (
    .DIN(WX690),
    .DIN_t(WX690_t),
    .SDIN(n6865),
    .SDIN_t(n6865_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6866),
    .Q_t(n6866_t),
    .QN(n6556),
    .QN_t(n6556_t)
  );


  sdffs1
  \DFF_54/Q_reg 
  (
    .DIN(WX688),
    .DIN_t(WX688_t),
    .SDIN(n6864),
    .SDIN_t(n6864_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6865),
    .Q_t(n6865_t),
    .QN(n6507),
    .QN_t(n6507_t)
  );


  sdffs1
  \DFF_53/Q_reg 
  (
    .DIN(WX686),
    .DIN_t(WX686_t),
    .SDIN(n6863),
    .SDIN_t(n6863_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6864),
    .Q_t(n6864_t),
    .QN(n6557),
    .QN_t(n6557_t)
  );


  sdffs1
  \DFF_52/Q_reg 
  (
    .DIN(WX684),
    .DIN_t(WX684_t),
    .SDIN(n6862),
    .SDIN_t(n6862_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6863),
    .Q_t(n6863_t),
    .QN(n6559),
    .QN_t(n6559_t)
  );


  sdffs1
  \DFF_51/Q_reg 
  (
    .DIN(WX682),
    .DIN_t(WX682_t),
    .SDIN(n6861),
    .SDIN_t(n6861_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6862),
    .Q_t(n6862_t),
    .QN(n6555),
    .QN_t(n6555_t)
  );


  sdffs1
  \DFF_50/Q_reg 
  (
    .DIN(WX680),
    .DIN_t(WX680_t),
    .SDIN(n6860),
    .SDIN_t(n6860_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6861),
    .Q_t(n6861_t),
    .QN(n6558),
    .QN_t(n6558_t)
  );


  sdffs1
  \DFF_49/Q_reg 
  (
    .DIN(WX678),
    .DIN_t(WX678_t),
    .SDIN(n6859),
    .SDIN_t(n6859_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6860),
    .Q_t(n6860_t),
    .QN(n6526),
    .QN_t(n6526_t)
  );


  sdffs1
  \DFF_48/Q_reg 
  (
    .DIN(WX676),
    .DIN_t(WX676_t),
    .SDIN(n6858),
    .SDIN_t(n6858_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6859),
    .Q_t(n6859_t),
    .QN(n6561),
    .QN_t(n6561_t)
  );


  sdffs1
  \DFF_47/Q_reg 
  (
    .DIN(WX674),
    .DIN_t(WX674_t),
    .SDIN(n6857),
    .SDIN_t(n6857_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6858),
    .Q_t(n6858_t),
    .QN(n6509),
    .QN_t(n6509_t)
  );


  sdffs1
  \DFF_46/Q_reg 
  (
    .DIN(WX672),
    .DIN_t(WX672_t),
    .SDIN(n6856),
    .SDIN_t(n6856_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6857),
    .Q_t(n6857_t),
    .QN(n6542),
    .QN_t(n6542_t)
  );


  sdffs1
  \DFF_45/Q_reg 
  (
    .DIN(WX670),
    .DIN_t(WX670_t),
    .SDIN(n6855),
    .SDIN_t(n6855_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6856),
    .Q_t(n6856_t),
    .QN(n6490),
    .QN_t(n6490_t)
  );


  sdffs1
  \DFF_44/Q_reg 
  (
    .DIN(WX668),
    .DIN_t(WX668_t),
    .SDIN(n6854),
    .SDIN_t(n6854_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6855),
    .Q_t(n6855_t),
    .QN(n6548),
    .QN_t(n6548_t)
  );


  sdffs1
  \DFF_43/Q_reg 
  (
    .DIN(WX666),
    .DIN_t(WX666_t),
    .SDIN(n6853),
    .SDIN_t(n6853_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6854),
    .Q_t(n6854_t),
    .QN(n6521),
    .QN_t(n6521_t)
  );


  sdffs1
  \DFF_42/Q_reg 
  (
    .DIN(WX664),
    .DIN_t(WX664_t),
    .SDIN(n6852),
    .SDIN_t(n6852_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6853),
    .Q_t(n6853_t),
    .QN(n6536),
    .QN_t(n6536_t)
  );


  sdffs1
  \DFF_41/Q_reg 
  (
    .DIN(WX662),
    .DIN_t(WX662_t),
    .SDIN(n6851),
    .SDIN_t(n6851_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6852),
    .Q_t(n6852_t),
    .QN(n6515),
    .QN_t(n6515_t)
  );


  sdffs1
  \DFF_40/Q_reg 
  (
    .DIN(WX660),
    .DIN_t(WX660_t),
    .SDIN(n6850),
    .SDIN_t(n6850_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6851),
    .Q_t(n6851_t),
    .QN(n6538),
    .QN_t(n6538_t)
  );


  sdffs1
  \DFF_39/Q_reg 
  (
    .DIN(WX658),
    .DIN_t(WX658_t),
    .SDIN(n6849),
    .SDIN_t(n6849_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6850),
    .Q_t(n6850_t),
    .QN(n6540),
    .QN_t(n6540_t)
  );


  sdffs1
  \DFF_38/Q_reg 
  (
    .DIN(WX656),
    .DIN_t(WX656_t),
    .SDIN(n6848),
    .SDIN_t(n6848_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6849),
    .Q_t(n6849_t),
    .QN(n6499),
    .QN_t(n6499_t)
  );


  sdffs1
  \DFF_37/Q_reg 
  (
    .DIN(WX654),
    .DIN_t(WX654_t),
    .SDIN(n6847),
    .SDIN_t(n6847_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6848),
    .Q_t(n6848_t),
    .QN(n6543),
    .QN_t(n6543_t)
  );


  sdffs1
  \DFF_36/Q_reg 
  (
    .DIN(WX652),
    .DIN_t(WX652_t),
    .SDIN(n6846),
    .SDIN_t(n6846_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6847),
    .Q_t(n6847_t),
    .QN(n6545),
    .QN_t(n6545_t)
  );


  sdffs1
  \DFF_35/Q_reg 
  (
    .DIN(WX650),
    .DIN_t(WX650_t),
    .SDIN(n6845),
    .SDIN_t(n6845_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6846),
    .Q_t(n6846_t),
    .QN(n6546),
    .QN_t(n6546_t)
  );


  sdffs1
  \DFF_34/Q_reg 
  (
    .DIN(WX648),
    .DIN_t(WX648_t),
    .SDIN(n6844),
    .SDIN_t(n6844_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6845),
    .Q_t(n6845_t),
    .QN(n6481),
    .QN_t(n6481_t)
  );


  sdffs1
  \DFF_33/Q_reg 
  (
    .DIN(WX646),
    .DIN_t(WX646_t),
    .SDIN(n6843),
    .SDIN_t(n6843_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6844),
    .Q_t(n6844_t),
    .QN(n6549),
    .QN_t(n6549_t)
  );


  sdffs1
  \DFF_32/Q_reg 
  (
    .DIN(WX644),
    .DIN_t(WX644_t),
    .SDIN(n6842),
    .SDIN_t(n6842_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6843),
    .Q_t(n6843_t),
    .QN(n6533),
    .QN_t(n6533_t)
  );


  sdffs1
  \DFF_31/Q_reg 
  (
    .DIN(WX546),
    .DIN_t(WX546_t),
    .SDIN(n6841),
    .SDIN_t(n6841_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6842),
    .Q_t(n6842_t),
    .QN(n6179),
    .QN_t(n6179_t)
  );


  sdffs1
  \DFF_30/Q_reg 
  (
    .DIN(WX544),
    .DIN_t(WX544_t),
    .SDIN(n6840),
    .SDIN_t(n6840_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6841),
    .Q_t(n6841_t),
    .QN(n6180),
    .QN_t(n6180_t)
  );


  sdffs1
  \DFF_29/Q_reg 
  (
    .DIN(WX542),
    .DIN_t(WX542_t),
    .SDIN(n6839),
    .SDIN_t(n6839_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6840),
    .Q_t(n6840_t),
    .QN(n6181),
    .QN_t(n6181_t)
  );


  sdffs1
  \DFF_28/Q_reg 
  (
    .DIN(WX540),
    .DIN_t(WX540_t),
    .SDIN(n6838),
    .SDIN_t(n6838_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6839),
    .Q_t(n6839_t),
    .QN(n6182),
    .QN_t(n6182_t)
  );


  sdffs1
  \DFF_27/Q_reg 
  (
    .DIN(WX538),
    .DIN_t(WX538_t),
    .SDIN(n6837),
    .SDIN_t(n6837_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6838),
    .Q_t(n6838_t),
    .QN(n6183),
    .QN_t(n6183_t)
  );


  sdffs1
  \DFF_26/Q_reg 
  (
    .DIN(WX536),
    .DIN_t(WX536_t),
    .SDIN(n6836),
    .SDIN_t(n6836_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6837),
    .Q_t(n6837_t),
    .QN(n6184),
    .QN_t(n6184_t)
  );


  sdffs1
  \DFF_25/Q_reg 
  (
    .DIN(WX534),
    .DIN_t(WX534_t),
    .SDIN(n6835),
    .SDIN_t(n6835_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6836),
    .Q_t(n6836_t),
    .QN(n6185),
    .QN_t(n6185_t)
  );


  sdffs1
  \DFF_24/Q_reg 
  (
    .DIN(WX532),
    .DIN_t(WX532_t),
    .SDIN(n6834),
    .SDIN_t(n6834_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6835),
    .Q_t(n6835_t),
    .QN(n6186),
    .QN_t(n6186_t)
  );


  sdffs1
  \DFF_23/Q_reg 
  (
    .DIN(WX530),
    .DIN_t(WX530_t),
    .SDIN(n6833),
    .SDIN_t(n6833_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6834),
    .Q_t(n6834_t),
    .QN(n6187),
    .QN_t(n6187_t)
  );


  sdffs1
  \DFF_22/Q_reg 
  (
    .DIN(WX528),
    .DIN_t(WX528_t),
    .SDIN(n6832),
    .SDIN_t(n6832_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6833),
    .Q_t(n6833_t),
    .QN(n6188),
    .QN_t(n6188_t)
  );


  sdffs1
  \DFF_21/Q_reg 
  (
    .DIN(WX526),
    .DIN_t(WX526_t),
    .SDIN(n6831),
    .SDIN_t(n6831_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6832),
    .Q_t(n6832_t),
    .QN(n6189),
    .QN_t(n6189_t)
  );


  sdffs1
  \DFF_20/Q_reg 
  (
    .DIN(WX524),
    .DIN_t(WX524_t),
    .SDIN(n6830),
    .SDIN_t(n6830_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6831),
    .Q_t(n6831_t),
    .QN(n6190),
    .QN_t(n6190_t)
  );


  sdffs1
  \DFF_19/Q_reg 
  (
    .DIN(WX522),
    .DIN_t(WX522_t),
    .SDIN(n6829),
    .SDIN_t(n6829_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6830),
    .Q_t(n6830_t),
    .QN(n6191),
    .QN_t(n6191_t)
  );


  sdffs1
  \DFF_18/Q_reg 
  (
    .DIN(WX520),
    .DIN_t(WX520_t),
    .SDIN(n6828),
    .SDIN_t(n6828_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6829),
    .Q_t(n6829_t),
    .QN(n6192),
    .QN_t(n6192_t)
  );


  sdffs1
  \DFF_17/Q_reg 
  (
    .DIN(WX518),
    .DIN_t(WX518_t),
    .SDIN(n6827),
    .SDIN_t(n6827_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6828),
    .Q_t(n6828_t),
    .QN(n6193),
    .QN_t(n6193_t)
  );


  sdffs1
  \DFF_16/Q_reg 
  (
    .DIN(WX516),
    .DIN_t(WX516_t),
    .SDIN(n6826),
    .SDIN_t(n6826_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6827),
    .Q_t(n6827_t),
    .QN(n6194),
    .QN_t(n6194_t)
  );


  sdffs1
  \DFF_15/Q_reg 
  (
    .DIN(WX514),
    .DIN_t(WX514_t),
    .SDIN(n6825),
    .SDIN_t(n6825_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6826),
    .Q_t(n6826_t),
    .QN(n6195),
    .QN_t(n6195_t)
  );


  sdffs1
  \DFF_14/Q_reg 
  (
    .DIN(WX512),
    .DIN_t(WX512_t),
    .SDIN(n6824),
    .SDIN_t(n6824_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6825),
    .Q_t(n6825_t),
    .QN(n6196),
    .QN_t(n6196_t)
  );


  sdffs1
  \DFF_13/Q_reg 
  (
    .DIN(WX510),
    .DIN_t(WX510_t),
    .SDIN(n6823),
    .SDIN_t(n6823_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6824),
    .Q_t(n6824_t),
    .QN(n6286),
    .QN_t(n6286_t)
  );


  sdffs1
  \DFF_12/Q_reg 
  (
    .DIN(WX508),
    .DIN_t(WX508_t),
    .SDIN(n6822),
    .SDIN_t(n6822_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6823),
    .Q_t(n6823_t),
    .QN(n6342),
    .QN_t(n6342_t)
  );


  sdffs1
  \DFF_11/Q_reg 
  (
    .DIN(WX506),
    .DIN_t(WX506_t),
    .SDIN(n6821),
    .SDIN_t(n6821_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6822),
    .Q_t(n6822_t),
    .QN(n6354),
    .QN_t(n6354_t)
  );


  sdffs1
  \DFF_10/Q_reg 
  (
    .DIN(WX504),
    .DIN_t(WX504_t),
    .SDIN(n6820),
    .SDIN_t(n6820_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6821),
    .Q_t(n6821_t),
    .QN(n6376),
    .QN_t(n6376_t)
  );


  sdffs1
  \DFF_9/Q_reg 
  (
    .DIN(WX502),
    .DIN_t(WX502_t),
    .SDIN(n6819),
    .SDIN_t(n6819_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6820),
    .Q_t(n6820_t),
    .QN(n6377),
    .QN_t(n6377_t)
  );


  sdffs1
  \DFF_8/Q_reg 
  (
    .DIN(WX500),
    .DIN_t(WX500_t),
    .SDIN(n6818),
    .SDIN_t(n6818_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6819),
    .Q_t(n6819_t),
    .QN(n6378),
    .QN_t(n6378_t)
  );


  sdffs1
  \DFF_7/Q_reg 
  (
    .DIN(WX498),
    .DIN_t(WX498_t),
    .SDIN(n6817),
    .SDIN_t(n6817_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6818),
    .Q_t(n6818_t),
    .QN(n6379),
    .QN_t(n6379_t)
  );


  sdffs1
  \DFF_6/Q_reg 
  (
    .DIN(WX496),
    .DIN_t(WX496_t),
    .SDIN(n6816),
    .SDIN_t(n6816_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6817),
    .Q_t(n6817_t),
    .QN(n6380),
    .QN_t(n6380_t)
  );


  sdffs1
  \DFF_5/Q_reg 
  (
    .DIN(WX494),
    .DIN_t(WX494_t),
    .SDIN(n6815),
    .SDIN_t(n6815_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6816),
    .Q_t(n6816_t),
    .QN(n6381),
    .QN_t(n6381_t)
  );


  sdffs1
  \DFF_4/Q_reg 
  (
    .DIN(WX492),
    .DIN_t(WX492_t),
    .SDIN(n6814),
    .SDIN_t(n6814_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6815),
    .Q_t(n6815_t),
    .QN(n6382),
    .QN_t(n6382_t)
  );


  sdffs1
  \DFF_3/Q_reg 
  (
    .DIN(WX490),
    .DIN_t(WX490_t),
    .SDIN(n6813),
    .SDIN_t(n6813_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6814),
    .Q_t(n6814_t),
    .QN(n6431),
    .QN_t(n6431_t)
  );


  sdffs1
  \DFF_2/Q_reg 
  (
    .DIN(WX488),
    .DIN_t(WX488_t),
    .SDIN(n6812),
    .SDIN_t(n6812_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6813),
    .Q_t(n6813_t),
    .QN(n6432),
    .QN_t(n6432_t)
  );


  sdffs1
  \DFF_1/Q_reg 
  (
    .DIN(WX486),
    .DIN_t(WX486_t),
    .SDIN(n6811),
    .SDIN_t(n6811_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6812),
    .Q_t(n6812_t),
    .QN(n6433),
    .QN_t(n6433_t)
  );


  sdffs1
  \DFF_0/Q_reg 
  (
    .DIN(WX484),
    .DIN_t(WX484_t),
    .SDIN(test_si),
    .SDIN_t(test_si_t),
    .SSEL(test_se),
    .SSEL_t(test_se_t),
    .CLK(CK),
    .CLK_t(CK_t),
    .Q(n6811),
    .Q_t(n6811_t),
    .QN(n6434),
    .QN_t(n6434_t)
  );


  nor4s1
  troj10_0U1
  (
    .DIN1(troj10_0n1),
    .DIN1_t(troj10_0n1_t),
    .DIN2(troj10_0n2),
    .DIN2_t(troj10_0n2_t),
    .DIN3(troj10_0n3),
    .DIN3_t(troj10_0n3_t),
    .DIN4(troj10_0n4),
    .DIN4_t(troj10_0n4_t),
    .Q(Trigger_en10_0),
    .Q_t(Trigger_en10_0_t)
  );


  nnd2s1
  troj10_0U2
  (
    .DIN1(n6564),
    .DIN1_t(n6564_t),
    .DIN2(n4549),
    .DIN2_t(n4549_t),
    .Q(troj10_0n4),
    .Q_t(troj10_0n4_t)
  );


  nnd2s1
  troj10_0U3
  (
    .DIN1(troj10_0n5),
    .DIN1_t(troj10_0n5_t),
    .DIN2(n4219),
    .DIN2_t(n4219_t),
    .Q(troj10_0n3),
    .Q_t(troj10_0n3_t)
  );


  and2s1
  troj10_0U4
  (
    .DIN1(n3359),
    .DIN1_t(n3359_t),
    .DIN2(n2954),
    .DIN2_t(n2954_t),
    .Q(troj10_0n5),
    .Q_t(troj10_0n5_t)
  );


  nnd2s1
  troj10_0U5
  (
    .DIN1(n2534),
    .DIN1_t(n2534_t),
    .DIN2(troj10_0n6),
    .DIN2_t(troj10_0n6_t),
    .Q(troj10_0n2),
    .Q_t(troj10_0n2_t)
  );


  i1s1
  troj10_0U6
  (
    .DIN(n1792),
    .DIN_t(n1792_t),
    .Q(troj10_0n6),
    .Q_t(troj10_0n6_t)
  );


  or3s1
  troj10_0U7
  (
    .DIN1(n2153),
    .DIN1_t(n2153_t),
    .DIN2(n1997),
    .DIN2_t(n1997_t),
    .DIN3(n1848),
    .DIN3_t(n1848_t),
    .Q(troj10_0n1),
    .Q_t(troj10_0n1_t)
  );


  xor2s1
  trojan10_0
  (
    .DIN1(tempn3869),
    .DIN1_t(tempn3869_t),
    .DIN2(Trigger_en10_0),
    .DIN2_t(Trigger_en10_0_t),
    .Q(n3869),
    .Q_t(n3869_t)
  );


  nor2s1
  troj10_1U1
  (
    .DIN1(troj10_1n1),
    .DIN1_t(troj10_1n1_t),
    .DIN2(troj10_1n2),
    .DIN2_t(troj10_1n2_t),
    .Q(Trigger_en10_1),
    .Q_t(Trigger_en10_1_t)
  );


  nnd4s1
  troj10_1U2
  (
    .DIN1(n4466),
    .DIN1_t(n4466_t),
    .DIN2(WX7011),
    .DIN2_t(WX7011_t),
    .DIN3(troj10_1n3),
    .DIN3_t(troj10_1n3_t),
    .DIN4(WX3882),
    .DIN4_t(WX3882_t),
    .Q(troj10_1n2),
    .Q_t(troj10_1n2_t)
  );


  nor2s1
  troj10_1U3
  (
    .DIN1(n1830),
    .DIN1_t(n1830_t),
    .DIN2(n1755),
    .DIN2_t(n1755_t),
    .Q(troj10_1n3),
    .Q_t(troj10_1n3_t)
  );


  or4s1
  troj10_1U4
  (
    .DIN1(n2579),
    .DIN1_t(n2579_t),
    .DIN2(n1958),
    .DIN2_t(n1958_t),
    .DIN3(n1931),
    .DIN3_t(n1931_t),
    .DIN4(troj10_1n4),
    .DIN4_t(troj10_1n4_t),
    .Q(troj10_1n1),
    .Q_t(troj10_1n1_t)
  );


  or3s1
  troj10_1U5
  (
    .DIN1(n3585),
    .DIN1_t(n3585_t),
    .DIN2(n3402),
    .DIN2_t(n3402_t),
    .DIN3(n3022),
    .DIN3_t(n3022_t),
    .Q(troj10_1n4),
    .Q_t(troj10_1n4_t)
  );


  xor2s1
  trojan10_1
  (
    .DIN1(tempn2493),
    .DIN1_t(tempn2493_t),
    .DIN2(Trigger_en10_1),
    .DIN2_t(Trigger_en10_1_t),
    .Q(n2493),
    .Q_t(n2493_t)
  );


endmodule

